VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO tt_um_JamesTimothyMeech_inverter
  CLASS BLOCK ;
  FOREIGN tt_um_JamesTimothyMeech_inverter ;
  ORIGIN 0.000 0.000 ;
  SIZE 161.000 BY 225.760 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 154.870 224.760 155.170 225.760 ;
    END
  END clk
  PIN ena
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 158.550 224.760 158.850 225.760 ;
    END
  END ena
  PIN rst_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 151.190 224.760 151.490 225.760 ;
    END
  END rst_n
  PIN ua[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 215.324997 ;
    PORT
      LAYER met4 ;
        RECT 156.560 0.000 157.160 1.000 ;
    END
  END ua[0]
  PIN ua[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 134.480 0.000 135.080 1.000 ;
    END
  END ua[1]
  PIN ua[2]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 112.400 0.000 113.000 1.000 ;
    END
  END ua[2]
  PIN ua[3]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 90.320 0.000 90.920 1.000 ;
    END
  END ua[3]
  PIN ua[4]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 5.800000 ;
    PORT
      LAYER met4 ;
        RECT 68.240 0.000 68.840 1.000 ;
    END
  END ua[4]
  PIN ua[5]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 20.000000 ;
    PORT
      LAYER met4 ;
        RECT 46.160 0.000 46.760 1.000 ;
    END
  END ua[5]
  PIN ua[6]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 24.080 0.000 24.680 1.000 ;
    END
  END ua[6]
  PIN ua[7]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 2.000 0.000 2.600 1.000 ;
    END
  END ua[7]
  PIN ui_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.675000 ;
    PORT
      LAYER met4 ;
        RECT 147.510 224.760 147.810 225.760 ;
    END
  END ui_in[0]
  PIN ui_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.675000 ;
    PORT
      LAYER met4 ;
        RECT 143.830 224.760 144.130 225.760 ;
    END
  END ui_in[1]
  PIN ui_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.675000 ;
    PORT
      LAYER met4 ;
        RECT 140.150 224.760 140.450 225.760 ;
    END
  END ui_in[2]
  PIN ui_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.675000 ;
    PORT
      LAYER met4 ;
        RECT 136.470 224.760 136.770 225.760 ;
    END
  END ui_in[3]
  PIN ui_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.675000 ;
    PORT
      LAYER met4 ;
        RECT 132.790 224.760 133.090 225.760 ;
    END
  END ui_in[4]
  PIN ui_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.675000 ;
    PORT
      LAYER met4 ;
        RECT 129.110 224.760 129.410 225.760 ;
    END
  END ui_in[5]
  PIN ui_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.675000 ;
    PORT
      LAYER met4 ;
        RECT 125.430 224.760 125.730 225.760 ;
    END
  END ui_in[6]
  PIN ui_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.675000 ;
    PORT
      LAYER met4 ;
        RECT 121.750 224.760 122.050 225.760 ;
    END
  END ui_in[7]
  PIN uio_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.675000 ;
    PORT
      LAYER met4 ;
        RECT 118.070 224.760 118.370 225.760 ;
    END
  END uio_in[0]
  PIN uio_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.675000 ;
    PORT
      LAYER met4 ;
        RECT 114.390 224.760 114.690 225.760 ;
    END
  END uio_in[1]
  PIN uio_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.675000 ;
    PORT
      LAYER met4 ;
        RECT 110.710 224.760 111.010 225.760 ;
    END
  END uio_in[2]
  PIN uio_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 107.030 224.760 107.330 225.760 ;
    END
  END uio_in[3]
  PIN uio_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 103.350 224.760 103.650 225.760 ;
    END
  END uio_in[4]
  PIN uio_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 99.670 224.760 99.970 225.760 ;
    END
  END uio_in[5]
  PIN uio_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 95.990 224.760 96.290 225.760 ;
    END
  END uio_in[6]
  PIN uio_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 92.310 224.760 92.610 225.760 ;
    END
  END uio_in[7]
  PIN uio_oe[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 152.991989 ;
    PORT
      LAYER met4 ;
        RECT 29.750 224.760 30.050 225.760 ;
    END
  END uio_oe[0]
  PIN uio_oe[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 152.991989 ;
    PORT
      LAYER met4 ;
        RECT 26.070 224.760 26.370 225.760 ;
    END
  END uio_oe[1]
  PIN uio_oe[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 152.991989 ;
    PORT
      LAYER met4 ;
        RECT 22.390 224.760 22.690 225.760 ;
    END
  END uio_oe[2]
  PIN uio_oe[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 152.991989 ;
    PORT
      LAYER met4 ;
        RECT 18.710 224.760 19.010 225.760 ;
    END
  END uio_oe[3]
  PIN uio_oe[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 152.991989 ;
    PORT
      LAYER met4 ;
        RECT 15.030 224.760 15.330 225.760 ;
    END
  END uio_oe[4]
  PIN uio_oe[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 152.991989 ;
    PORT
      LAYER met4 ;
        RECT 11.350 224.760 11.650 225.760 ;
    END
  END uio_oe[5]
  PIN uio_oe[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 152.991989 ;
    PORT
      LAYER met4 ;
        RECT 7.670 224.760 7.970 225.760 ;
    END
  END uio_oe[6]
  PIN uio_oe[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 152.991989 ;
    PORT
      LAYER met4 ;
        RECT 3.990 224.760 4.290 225.760 ;
    END
  END uio_oe[7]
  PIN uio_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 152.991989 ;
    PORT
      LAYER met4 ;
        RECT 59.190 224.760 59.490 225.760 ;
    END
  END uio_out[0]
  PIN uio_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 152.991989 ;
    PORT
      LAYER met4 ;
        RECT 55.510 224.760 55.810 225.760 ;
    END
  END uio_out[1]
  PIN uio_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 152.991989 ;
    PORT
      LAYER met4 ;
        RECT 51.830 224.760 52.130 225.760 ;
    END
  END uio_out[2]
  PIN uio_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 152.991989 ;
    PORT
      LAYER met4 ;
        RECT 48.150 224.760 48.450 225.760 ;
    END
  END uio_out[3]
  PIN uio_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 152.991989 ;
    PORT
      LAYER met4 ;
        RECT 44.470 224.760 44.770 225.760 ;
    END
  END uio_out[4]
  PIN uio_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 152.991989 ;
    PORT
      LAYER met4 ;
        RECT 40.790 224.760 41.090 225.760 ;
    END
  END uio_out[5]
  PIN uio_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 152.991989 ;
    PORT
      LAYER met4 ;
        RECT 37.110 224.760 37.410 225.760 ;
    END
  END uio_out[6]
  PIN uio_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 152.991989 ;
    PORT
      LAYER met4 ;
        RECT 33.430 224.760 33.730 225.760 ;
    END
  END uio_out[7]
  PIN uo_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 152.991989 ;
    PORT
      LAYER met4 ;
        RECT 88.630 224.760 88.930 225.760 ;
    END
  END uo_out[0]
  PIN uo_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 152.991989 ;
    PORT
      LAYER met4 ;
        RECT 84.950 224.760 85.250 225.760 ;
    END
  END uo_out[1]
  PIN uo_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 152.991989 ;
    PORT
      LAYER met4 ;
        RECT 81.270 224.760 81.570 225.760 ;
    END
  END uo_out[2]
  PIN uo_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 152.991989 ;
    PORT
      LAYER met4 ;
        RECT 77.590 224.760 77.890 225.760 ;
    END
  END uo_out[3]
  PIN uo_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 152.991989 ;
    PORT
      LAYER met4 ;
        RECT 73.910 224.760 74.210 225.760 ;
    END
  END uo_out[4]
  PIN uo_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 152.991989 ;
    PORT
      LAYER met4 ;
        RECT 70.230 224.760 70.530 225.760 ;
    END
  END uo_out[5]
  PIN uo_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 152.991989 ;
    PORT
      LAYER met4 ;
        RECT 66.550 224.760 66.850 225.760 ;
    END
  END uo_out[6]
  PIN uo_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 152.991989 ;
    PORT
      LAYER met4 ;
        RECT 62.870 224.760 63.170 225.760 ;
    END
  END uo_out[7]
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1.000 5.000 2.500 220.760 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 49.000 5.000 50.500 220.760 ;
    END
  END VGND
  OBS
      LAYER pwell ;
        RECT 60.790 199.580 62.800 199.780 ;
        RECT 59.490 198.200 62.800 199.580 ;
        RECT 60.790 183.800 62.800 198.200 ;
      LAYER nwell ;
        RECT 64.540 183.890 71.230 199.000 ;
        RECT 72.510 195.210 76.200 199.940 ;
      LAYER pwell ;
        RECT 85.530 199.500 87.540 199.700 ;
        RECT 76.400 195.730 80.000 199.420 ;
        RECT 84.230 198.120 87.540 199.500 ;
        RECT 73.000 187.830 79.600 193.980 ;
        RECT 85.530 183.720 87.540 198.120 ;
      LAYER nwell ;
        RECT 89.280 183.810 95.970 198.920 ;
        RECT 97.250 195.130 100.940 199.860 ;
      LAYER pwell ;
        RECT 108.780 199.490 110.790 199.690 ;
        RECT 101.140 195.650 104.740 199.340 ;
        RECT 107.480 198.110 110.790 199.490 ;
        RECT 97.740 187.750 104.340 193.900 ;
        RECT 108.780 183.710 110.790 198.110 ;
      LAYER nwell ;
        RECT 112.530 183.800 119.220 198.910 ;
        RECT 120.500 195.120 124.190 199.850 ;
      LAYER pwell ;
        RECT 132.410 199.480 134.420 199.680 ;
        RECT 124.390 195.640 127.990 199.330 ;
        RECT 131.110 198.100 134.420 199.480 ;
        RECT 120.990 187.740 127.590 193.890 ;
        RECT 132.410 183.700 134.420 198.100 ;
      LAYER nwell ;
        RECT 136.160 183.790 142.850 198.900 ;
        RECT 144.130 195.110 147.820 199.840 ;
      LAYER pwell ;
        RECT 148.020 195.630 151.620 199.320 ;
        RECT 144.620 187.730 151.220 193.880 ;
        RECT 60.680 173.490 62.690 173.690 ;
        RECT 59.380 172.110 62.690 173.490 ;
        RECT 60.680 157.710 62.690 172.110 ;
      LAYER nwell ;
        RECT 64.430 157.800 71.120 172.910 ;
        RECT 72.400 169.120 76.090 173.850 ;
      LAYER pwell ;
        RECT 83.860 173.400 85.870 173.600 ;
        RECT 76.290 169.640 79.890 173.330 ;
        RECT 82.560 172.020 85.870 173.400 ;
        RECT 72.890 161.740 79.490 167.890 ;
        RECT 83.860 157.620 85.870 172.020 ;
      LAYER nwell ;
        RECT 87.610 157.710 94.300 172.820 ;
        RECT 95.580 169.030 99.270 173.760 ;
      LAYER pwell ;
        RECT 106.760 173.600 108.770 173.800 ;
        RECT 99.470 169.550 103.070 173.240 ;
        RECT 105.460 172.220 108.770 173.600 ;
        RECT 96.070 161.650 102.670 167.800 ;
        RECT 106.760 157.820 108.770 172.220 ;
      LAYER nwell ;
        RECT 110.510 157.910 117.200 173.020 ;
        RECT 118.480 169.230 122.170 173.960 ;
      LAYER pwell ;
        RECT 129.860 173.710 131.870 173.910 ;
        RECT 122.370 169.750 125.970 173.440 ;
        RECT 128.560 172.330 131.870 173.710 ;
        RECT 118.970 161.850 125.570 168.000 ;
        RECT 129.860 157.930 131.870 172.330 ;
      LAYER nwell ;
        RECT 133.610 158.020 140.300 173.130 ;
        RECT 141.580 169.340 145.270 174.070 ;
      LAYER pwell ;
        RECT 145.470 169.860 149.070 173.550 ;
        RECT 142.070 161.960 148.670 168.110 ;
        RECT 84.070 147.760 86.080 147.960 ;
        RECT 82.770 146.380 86.080 147.760 ;
        RECT 84.070 131.980 86.080 146.380 ;
      LAYER nwell ;
        RECT 87.820 132.070 94.510 147.180 ;
        RECT 95.790 143.390 99.480 148.120 ;
      LAYER pwell ;
        RECT 107.100 147.910 109.110 148.110 ;
        RECT 99.680 143.910 103.280 147.600 ;
        RECT 105.800 146.530 109.110 147.910 ;
        RECT 96.280 136.010 102.880 142.160 ;
        RECT 107.100 132.130 109.110 146.530 ;
      LAYER nwell ;
        RECT 110.850 132.220 117.540 147.330 ;
        RECT 118.820 143.540 122.510 148.270 ;
      LAYER pwell ;
        RECT 130.110 147.990 132.120 148.190 ;
        RECT 122.710 144.060 126.310 147.750 ;
        RECT 128.810 146.610 132.120 147.990 ;
        RECT 119.310 136.160 125.910 142.310 ;
        RECT 130.110 132.210 132.120 146.610 ;
      LAYER nwell ;
        RECT 133.860 132.300 140.550 147.410 ;
        RECT 141.830 143.620 145.520 148.350 ;
      LAYER pwell ;
        RECT 145.720 144.140 149.320 147.830 ;
        RECT 142.320 136.240 148.920 142.390 ;
      LAYER nwell ;
        RECT 57.550 22.720 60.510 34.910 ;
      LAYER pwell ;
        RECT 57.500 16.280 60.460 17.430 ;
        RECT 57.500 6.480 60.520 16.280 ;
        RECT 57.500 5.330 60.460 6.480 ;
      LAYER li1 ;
        RECT 61.450 199.600 62.140 199.610 ;
        RECT 60.970 199.430 62.620 199.600 ;
        RECT 72.690 199.590 76.020 199.760 ;
        RECT 72.690 199.510 72.860 199.590 ;
        RECT 60.970 184.150 61.140 199.430 ;
        RECT 61.620 196.790 61.970 198.950 ;
        RECT 61.620 184.630 61.970 186.790 ;
        RECT 62.450 184.150 62.620 199.430 ;
        RECT 70.880 198.820 72.860 199.510 ;
        RECT 60.970 183.980 62.620 184.150 ;
        RECT 64.720 198.650 72.860 198.820 ;
        RECT 64.720 184.240 64.890 198.650 ;
        RECT 65.615 198.080 70.155 198.250 ;
        RECT 65.230 197.670 65.400 198.020 ;
        RECT 70.370 197.670 70.540 198.020 ;
        RECT 70.880 197.660 72.860 198.650 ;
        RECT 73.195 198.215 73.375 199.035 ;
        RECT 73.585 199.020 75.125 199.190 ;
        RECT 73.585 198.540 75.125 198.710 ;
        RECT 73.585 198.060 75.125 198.230 ;
        RECT 75.335 198.215 75.515 199.035 ;
        RECT 75.850 197.660 76.020 199.590 ;
        RECT 86.190 199.520 86.880 199.530 ;
        RECT 79.640 199.240 81.300 199.510 ;
        RECT 65.615 197.440 70.155 197.610 ;
        RECT 70.880 197.490 76.020 197.660 ;
        RECT 65.230 197.030 65.400 197.380 ;
        RECT 70.370 197.030 70.540 197.380 ;
        RECT 65.615 196.800 70.155 196.970 ;
        RECT 65.230 196.390 65.400 196.740 ;
        RECT 70.370 196.390 70.540 196.740 ;
        RECT 65.615 196.160 70.155 196.330 ;
        RECT 65.230 195.750 65.400 196.100 ;
        RECT 70.370 195.750 70.540 196.100 ;
        RECT 65.615 195.520 70.155 195.690 ;
        RECT 70.880 195.560 72.860 197.490 ;
        RECT 73.195 196.115 73.375 196.935 ;
        RECT 73.585 196.920 75.125 197.090 ;
        RECT 73.585 196.440 75.125 196.610 ;
        RECT 73.585 195.960 75.125 196.130 ;
        RECT 75.335 196.115 75.515 196.935 ;
        RECT 75.850 195.560 76.020 197.490 ;
        RECT 76.580 199.070 81.300 199.240 ;
        RECT 76.580 197.660 76.750 199.070 ;
        RECT 77.090 198.200 77.260 198.530 ;
        RECT 77.430 198.500 78.970 198.670 ;
        RECT 77.430 198.060 78.970 198.230 ;
        RECT 79.140 198.200 79.310 198.530 ;
        RECT 79.640 197.660 81.300 199.070 ;
        RECT 76.580 197.490 81.300 197.660 ;
        RECT 76.580 196.080 76.750 197.490 ;
        RECT 77.090 196.620 77.260 196.950 ;
        RECT 77.430 196.920 78.970 197.090 ;
        RECT 77.430 196.480 78.970 196.650 ;
        RECT 79.140 196.620 79.310 196.950 ;
        RECT 79.640 196.080 81.300 197.490 ;
        RECT 76.580 195.910 81.300 196.080 ;
        RECT 65.230 195.110 65.400 195.460 ;
        RECT 70.370 195.110 70.540 195.460 ;
        RECT 70.880 195.390 76.020 195.560 ;
        RECT 65.615 194.880 70.155 195.050 ;
        RECT 65.230 194.470 65.400 194.820 ;
        RECT 70.370 194.470 70.540 194.820 ;
        RECT 65.615 194.240 70.155 194.410 ;
        RECT 65.230 193.830 65.400 194.180 ;
        RECT 70.370 193.830 70.540 194.180 ;
        RECT 65.615 193.600 70.155 193.770 ;
        RECT 65.230 193.190 65.400 193.540 ;
        RECT 70.370 193.190 70.540 193.540 ;
        RECT 65.615 192.960 70.155 193.130 ;
        RECT 65.230 192.550 65.400 192.900 ;
        RECT 70.370 192.550 70.540 192.900 ;
        RECT 65.615 192.320 70.155 192.490 ;
        RECT 65.230 191.910 65.400 192.260 ;
        RECT 70.370 191.910 70.540 192.260 ;
        RECT 65.615 191.680 70.155 191.850 ;
        RECT 65.230 191.270 65.400 191.620 ;
        RECT 70.370 191.270 70.540 191.620 ;
        RECT 65.615 191.040 70.155 191.210 ;
        RECT 65.230 190.630 65.400 190.980 ;
        RECT 70.370 190.630 70.540 190.980 ;
        RECT 65.615 190.400 70.155 190.570 ;
        RECT 65.230 189.990 65.400 190.340 ;
        RECT 70.370 189.990 70.540 190.340 ;
        RECT 65.615 189.760 70.155 189.930 ;
        RECT 65.230 189.350 65.400 189.700 ;
        RECT 70.370 189.350 70.540 189.700 ;
        RECT 65.615 189.120 70.155 189.290 ;
        RECT 65.230 188.710 65.400 189.060 ;
        RECT 70.370 188.710 70.540 189.060 ;
        RECT 65.615 188.480 70.155 188.650 ;
        RECT 65.230 188.070 65.400 188.420 ;
        RECT 70.370 188.070 70.540 188.420 ;
        RECT 65.615 187.840 70.155 188.010 ;
        RECT 65.230 187.430 65.400 187.780 ;
        RECT 70.370 187.430 70.540 187.780 ;
        RECT 65.615 187.200 70.155 187.370 ;
        RECT 65.230 186.790 65.400 187.140 ;
        RECT 70.370 186.790 70.540 187.140 ;
        RECT 65.615 186.560 70.155 186.730 ;
        RECT 65.230 186.150 65.400 186.500 ;
        RECT 70.370 186.150 70.540 186.500 ;
        RECT 65.615 185.920 70.155 186.090 ;
        RECT 65.230 185.510 65.400 185.860 ;
        RECT 70.370 185.510 70.540 185.860 ;
        RECT 65.615 185.280 70.155 185.450 ;
        RECT 65.230 184.870 65.400 185.220 ;
        RECT 70.370 184.870 70.540 185.220 ;
        RECT 65.615 184.640 70.155 184.810 ;
        RECT 70.880 184.240 72.500 195.390 ;
        RECT 79.640 193.800 81.300 195.910 ;
        RECT 73.180 193.630 81.300 193.800 ;
        RECT 73.180 188.180 73.350 193.630 ;
        RECT 74.030 193.060 78.570 193.230 ;
        RECT 73.690 192.650 73.860 193.000 ;
        RECT 78.740 192.650 78.910 193.000 ;
        RECT 74.030 192.420 78.570 192.590 ;
        RECT 73.690 192.010 73.860 192.360 ;
        RECT 78.740 192.010 78.910 192.360 ;
        RECT 74.030 191.780 78.570 191.950 ;
        RECT 73.690 191.370 73.860 191.720 ;
        RECT 78.740 191.370 78.910 191.720 ;
        RECT 74.030 191.140 78.570 191.310 ;
        RECT 73.690 190.730 73.860 191.080 ;
        RECT 78.740 190.730 78.910 191.080 ;
        RECT 74.030 190.500 78.570 190.670 ;
        RECT 73.690 190.090 73.860 190.440 ;
        RECT 78.740 190.090 78.910 190.440 ;
        RECT 74.030 189.860 78.570 190.030 ;
        RECT 73.690 189.450 73.860 189.800 ;
        RECT 78.740 189.450 78.910 189.800 ;
        RECT 74.030 189.220 78.570 189.390 ;
        RECT 73.690 188.810 73.860 189.160 ;
        RECT 78.740 188.810 78.910 189.160 ;
        RECT 74.030 188.580 78.570 188.750 ;
        RECT 79.250 188.180 81.300 193.630 ;
        RECT 73.180 188.010 81.300 188.180 ;
        RECT 64.720 184.070 72.500 184.240 ;
        RECT 70.880 182.310 72.500 184.070 ;
        RECT 80.100 182.310 81.300 188.010 ;
        RECT 85.710 199.350 87.360 199.520 ;
        RECT 97.430 199.510 100.760 199.680 ;
        RECT 109.440 199.510 110.130 199.520 ;
        RECT 97.430 199.430 97.600 199.510 ;
        RECT 85.710 184.070 85.880 199.350 ;
        RECT 86.360 196.710 86.710 198.870 ;
        RECT 86.360 184.550 86.710 186.710 ;
        RECT 87.190 184.070 87.360 199.350 ;
        RECT 95.620 198.740 97.600 199.430 ;
        RECT 85.710 183.900 87.360 184.070 ;
        RECT 89.460 198.570 97.600 198.740 ;
        RECT 89.460 184.160 89.630 198.570 ;
        RECT 90.355 198.000 94.895 198.170 ;
        RECT 89.970 197.590 90.140 197.940 ;
        RECT 95.110 197.590 95.280 197.940 ;
        RECT 95.620 197.580 97.600 198.570 ;
        RECT 97.935 198.135 98.115 198.955 ;
        RECT 98.325 198.940 99.865 199.110 ;
        RECT 98.325 198.460 99.865 198.630 ;
        RECT 98.325 197.980 99.865 198.150 ;
        RECT 100.075 198.135 100.255 198.955 ;
        RECT 100.590 197.580 100.760 199.510 ;
        RECT 104.380 199.160 106.040 199.430 ;
        RECT 90.355 197.360 94.895 197.530 ;
        RECT 95.620 197.410 100.760 197.580 ;
        RECT 89.970 196.950 90.140 197.300 ;
        RECT 95.110 196.950 95.280 197.300 ;
        RECT 90.355 196.720 94.895 196.890 ;
        RECT 89.970 196.310 90.140 196.660 ;
        RECT 95.110 196.310 95.280 196.660 ;
        RECT 90.355 196.080 94.895 196.250 ;
        RECT 89.970 195.670 90.140 196.020 ;
        RECT 95.110 195.670 95.280 196.020 ;
        RECT 90.355 195.440 94.895 195.610 ;
        RECT 95.620 195.480 97.600 197.410 ;
        RECT 97.935 196.035 98.115 196.855 ;
        RECT 98.325 196.840 99.865 197.010 ;
        RECT 98.325 196.360 99.865 196.530 ;
        RECT 98.325 195.880 99.865 196.050 ;
        RECT 100.075 196.035 100.255 196.855 ;
        RECT 100.590 195.480 100.760 197.410 ;
        RECT 101.320 198.990 106.040 199.160 ;
        RECT 101.320 197.580 101.490 198.990 ;
        RECT 101.830 198.120 102.000 198.450 ;
        RECT 102.170 198.420 103.710 198.590 ;
        RECT 102.170 197.980 103.710 198.150 ;
        RECT 103.880 198.120 104.050 198.450 ;
        RECT 104.380 197.580 106.040 198.990 ;
        RECT 101.320 197.410 106.040 197.580 ;
        RECT 101.320 196.000 101.490 197.410 ;
        RECT 101.830 196.540 102.000 196.870 ;
        RECT 102.170 196.840 103.710 197.010 ;
        RECT 102.170 196.400 103.710 196.570 ;
        RECT 103.880 196.540 104.050 196.870 ;
        RECT 104.380 196.000 106.040 197.410 ;
        RECT 101.320 195.830 106.040 196.000 ;
        RECT 89.970 195.030 90.140 195.380 ;
        RECT 95.110 195.030 95.280 195.380 ;
        RECT 95.620 195.310 100.760 195.480 ;
        RECT 90.355 194.800 94.895 194.970 ;
        RECT 89.970 194.390 90.140 194.740 ;
        RECT 95.110 194.390 95.280 194.740 ;
        RECT 90.355 194.160 94.895 194.330 ;
        RECT 89.970 193.750 90.140 194.100 ;
        RECT 95.110 193.750 95.280 194.100 ;
        RECT 90.355 193.520 94.895 193.690 ;
        RECT 89.970 193.110 90.140 193.460 ;
        RECT 95.110 193.110 95.280 193.460 ;
        RECT 90.355 192.880 94.895 193.050 ;
        RECT 89.970 192.470 90.140 192.820 ;
        RECT 95.110 192.470 95.280 192.820 ;
        RECT 90.355 192.240 94.895 192.410 ;
        RECT 89.970 191.830 90.140 192.180 ;
        RECT 95.110 191.830 95.280 192.180 ;
        RECT 90.355 191.600 94.895 191.770 ;
        RECT 89.970 191.190 90.140 191.540 ;
        RECT 95.110 191.190 95.280 191.540 ;
        RECT 90.355 190.960 94.895 191.130 ;
        RECT 89.970 190.550 90.140 190.900 ;
        RECT 95.110 190.550 95.280 190.900 ;
        RECT 90.355 190.320 94.895 190.490 ;
        RECT 89.970 189.910 90.140 190.260 ;
        RECT 95.110 189.910 95.280 190.260 ;
        RECT 90.355 189.680 94.895 189.850 ;
        RECT 89.970 189.270 90.140 189.620 ;
        RECT 95.110 189.270 95.280 189.620 ;
        RECT 90.355 189.040 94.895 189.210 ;
        RECT 89.970 188.630 90.140 188.980 ;
        RECT 95.110 188.630 95.280 188.980 ;
        RECT 90.355 188.400 94.895 188.570 ;
        RECT 89.970 187.990 90.140 188.340 ;
        RECT 95.110 187.990 95.280 188.340 ;
        RECT 90.355 187.760 94.895 187.930 ;
        RECT 89.970 187.350 90.140 187.700 ;
        RECT 95.110 187.350 95.280 187.700 ;
        RECT 90.355 187.120 94.895 187.290 ;
        RECT 89.970 186.710 90.140 187.060 ;
        RECT 95.110 186.710 95.280 187.060 ;
        RECT 90.355 186.480 94.895 186.650 ;
        RECT 89.970 186.070 90.140 186.420 ;
        RECT 95.110 186.070 95.280 186.420 ;
        RECT 90.355 185.840 94.895 186.010 ;
        RECT 89.970 185.430 90.140 185.780 ;
        RECT 95.110 185.430 95.280 185.780 ;
        RECT 90.355 185.200 94.895 185.370 ;
        RECT 89.970 184.790 90.140 185.140 ;
        RECT 95.110 184.790 95.280 185.140 ;
        RECT 90.355 184.560 94.895 184.730 ;
        RECT 95.620 184.160 97.240 195.310 ;
        RECT 104.380 193.720 106.040 195.830 ;
        RECT 97.920 193.550 106.040 193.720 ;
        RECT 97.920 188.100 98.090 193.550 ;
        RECT 98.770 192.980 103.310 193.150 ;
        RECT 98.430 192.570 98.600 192.920 ;
        RECT 103.480 192.570 103.650 192.920 ;
        RECT 98.770 192.340 103.310 192.510 ;
        RECT 98.430 191.930 98.600 192.280 ;
        RECT 103.480 191.930 103.650 192.280 ;
        RECT 98.770 191.700 103.310 191.870 ;
        RECT 98.430 191.290 98.600 191.640 ;
        RECT 103.480 191.290 103.650 191.640 ;
        RECT 98.770 191.060 103.310 191.230 ;
        RECT 98.430 190.650 98.600 191.000 ;
        RECT 103.480 190.650 103.650 191.000 ;
        RECT 98.770 190.420 103.310 190.590 ;
        RECT 98.430 190.010 98.600 190.360 ;
        RECT 103.480 190.010 103.650 190.360 ;
        RECT 98.770 189.780 103.310 189.950 ;
        RECT 98.430 189.370 98.600 189.720 ;
        RECT 103.480 189.370 103.650 189.720 ;
        RECT 98.770 189.140 103.310 189.310 ;
        RECT 98.430 188.730 98.600 189.080 ;
        RECT 103.480 188.730 103.650 189.080 ;
        RECT 98.770 188.500 103.310 188.670 ;
        RECT 103.990 188.100 106.040 193.550 ;
        RECT 97.920 187.930 106.040 188.100 ;
        RECT 89.460 183.990 97.240 184.160 ;
        RECT 95.620 182.230 97.240 183.990 ;
        RECT 104.840 182.230 106.040 187.930 ;
        RECT 108.960 199.340 110.610 199.510 ;
        RECT 120.680 199.500 124.010 199.670 ;
        RECT 133.070 199.500 133.760 199.510 ;
        RECT 120.680 199.420 120.850 199.500 ;
        RECT 108.960 184.060 109.130 199.340 ;
        RECT 109.610 196.700 109.960 198.860 ;
        RECT 109.610 184.540 109.960 186.700 ;
        RECT 110.440 184.060 110.610 199.340 ;
        RECT 118.870 198.730 120.850 199.420 ;
        RECT 108.960 183.890 110.610 184.060 ;
        RECT 112.710 198.560 120.850 198.730 ;
        RECT 112.710 184.150 112.880 198.560 ;
        RECT 113.605 197.990 118.145 198.160 ;
        RECT 113.220 197.580 113.390 197.930 ;
        RECT 118.360 197.580 118.530 197.930 ;
        RECT 118.870 197.570 120.850 198.560 ;
        RECT 121.185 198.125 121.365 198.945 ;
        RECT 121.575 198.930 123.115 199.100 ;
        RECT 121.575 198.450 123.115 198.620 ;
        RECT 121.575 197.970 123.115 198.140 ;
        RECT 123.325 198.125 123.505 198.945 ;
        RECT 123.840 197.570 124.010 199.500 ;
        RECT 127.630 199.150 129.290 199.420 ;
        RECT 113.605 197.350 118.145 197.520 ;
        RECT 118.870 197.400 124.010 197.570 ;
        RECT 113.220 196.940 113.390 197.290 ;
        RECT 118.360 196.940 118.530 197.290 ;
        RECT 113.605 196.710 118.145 196.880 ;
        RECT 113.220 196.300 113.390 196.650 ;
        RECT 118.360 196.300 118.530 196.650 ;
        RECT 113.605 196.070 118.145 196.240 ;
        RECT 113.220 195.660 113.390 196.010 ;
        RECT 118.360 195.660 118.530 196.010 ;
        RECT 113.605 195.430 118.145 195.600 ;
        RECT 118.870 195.470 120.850 197.400 ;
        RECT 121.185 196.025 121.365 196.845 ;
        RECT 121.575 196.830 123.115 197.000 ;
        RECT 121.575 196.350 123.115 196.520 ;
        RECT 121.575 195.870 123.115 196.040 ;
        RECT 123.325 196.025 123.505 196.845 ;
        RECT 123.840 195.470 124.010 197.400 ;
        RECT 124.570 198.980 129.290 199.150 ;
        RECT 124.570 197.570 124.740 198.980 ;
        RECT 125.080 198.110 125.250 198.440 ;
        RECT 125.420 198.410 126.960 198.580 ;
        RECT 125.420 197.970 126.960 198.140 ;
        RECT 127.130 198.110 127.300 198.440 ;
        RECT 127.630 197.570 129.290 198.980 ;
        RECT 124.570 197.400 129.290 197.570 ;
        RECT 124.570 195.990 124.740 197.400 ;
        RECT 125.080 196.530 125.250 196.860 ;
        RECT 125.420 196.830 126.960 197.000 ;
        RECT 125.420 196.390 126.960 196.560 ;
        RECT 127.130 196.530 127.300 196.860 ;
        RECT 127.630 195.990 129.290 197.400 ;
        RECT 124.570 195.820 129.290 195.990 ;
        RECT 113.220 195.020 113.390 195.370 ;
        RECT 118.360 195.020 118.530 195.370 ;
        RECT 118.870 195.300 124.010 195.470 ;
        RECT 113.605 194.790 118.145 194.960 ;
        RECT 113.220 194.380 113.390 194.730 ;
        RECT 118.360 194.380 118.530 194.730 ;
        RECT 113.605 194.150 118.145 194.320 ;
        RECT 113.220 193.740 113.390 194.090 ;
        RECT 118.360 193.740 118.530 194.090 ;
        RECT 113.605 193.510 118.145 193.680 ;
        RECT 113.220 193.100 113.390 193.450 ;
        RECT 118.360 193.100 118.530 193.450 ;
        RECT 113.605 192.870 118.145 193.040 ;
        RECT 113.220 192.460 113.390 192.810 ;
        RECT 118.360 192.460 118.530 192.810 ;
        RECT 113.605 192.230 118.145 192.400 ;
        RECT 113.220 191.820 113.390 192.170 ;
        RECT 118.360 191.820 118.530 192.170 ;
        RECT 113.605 191.590 118.145 191.760 ;
        RECT 113.220 191.180 113.390 191.530 ;
        RECT 118.360 191.180 118.530 191.530 ;
        RECT 113.605 190.950 118.145 191.120 ;
        RECT 113.220 190.540 113.390 190.890 ;
        RECT 118.360 190.540 118.530 190.890 ;
        RECT 113.605 190.310 118.145 190.480 ;
        RECT 113.220 189.900 113.390 190.250 ;
        RECT 118.360 189.900 118.530 190.250 ;
        RECT 113.605 189.670 118.145 189.840 ;
        RECT 113.220 189.260 113.390 189.610 ;
        RECT 118.360 189.260 118.530 189.610 ;
        RECT 113.605 189.030 118.145 189.200 ;
        RECT 113.220 188.620 113.390 188.970 ;
        RECT 118.360 188.620 118.530 188.970 ;
        RECT 113.605 188.390 118.145 188.560 ;
        RECT 113.220 187.980 113.390 188.330 ;
        RECT 118.360 187.980 118.530 188.330 ;
        RECT 113.605 187.750 118.145 187.920 ;
        RECT 113.220 187.340 113.390 187.690 ;
        RECT 118.360 187.340 118.530 187.690 ;
        RECT 113.605 187.110 118.145 187.280 ;
        RECT 113.220 186.700 113.390 187.050 ;
        RECT 118.360 186.700 118.530 187.050 ;
        RECT 113.605 186.470 118.145 186.640 ;
        RECT 113.220 186.060 113.390 186.410 ;
        RECT 118.360 186.060 118.530 186.410 ;
        RECT 113.605 185.830 118.145 186.000 ;
        RECT 113.220 185.420 113.390 185.770 ;
        RECT 118.360 185.420 118.530 185.770 ;
        RECT 113.605 185.190 118.145 185.360 ;
        RECT 113.220 184.780 113.390 185.130 ;
        RECT 118.360 184.780 118.530 185.130 ;
        RECT 113.605 184.550 118.145 184.720 ;
        RECT 118.870 184.150 120.490 195.300 ;
        RECT 127.630 193.710 129.290 195.820 ;
        RECT 121.170 193.540 129.290 193.710 ;
        RECT 121.170 188.090 121.340 193.540 ;
        RECT 122.020 192.970 126.560 193.140 ;
        RECT 121.680 192.560 121.850 192.910 ;
        RECT 126.730 192.560 126.900 192.910 ;
        RECT 122.020 192.330 126.560 192.500 ;
        RECT 121.680 191.920 121.850 192.270 ;
        RECT 126.730 191.920 126.900 192.270 ;
        RECT 122.020 191.690 126.560 191.860 ;
        RECT 121.680 191.280 121.850 191.630 ;
        RECT 126.730 191.280 126.900 191.630 ;
        RECT 122.020 191.050 126.560 191.220 ;
        RECT 121.680 190.640 121.850 190.990 ;
        RECT 126.730 190.640 126.900 190.990 ;
        RECT 122.020 190.410 126.560 190.580 ;
        RECT 121.680 190.000 121.850 190.350 ;
        RECT 126.730 190.000 126.900 190.350 ;
        RECT 122.020 189.770 126.560 189.940 ;
        RECT 121.680 189.360 121.850 189.710 ;
        RECT 126.730 189.360 126.900 189.710 ;
        RECT 122.020 189.130 126.560 189.300 ;
        RECT 121.680 188.720 121.850 189.070 ;
        RECT 126.730 188.720 126.900 189.070 ;
        RECT 122.020 188.490 126.560 188.660 ;
        RECT 127.240 188.090 129.290 193.540 ;
        RECT 121.170 187.920 129.290 188.090 ;
        RECT 112.710 183.980 120.490 184.150 ;
        RECT 118.870 182.220 120.490 183.980 ;
        RECT 128.090 182.220 129.290 187.920 ;
        RECT 132.590 199.330 134.240 199.500 ;
        RECT 144.310 199.490 147.640 199.660 ;
        RECT 144.310 199.410 144.480 199.490 ;
        RECT 132.590 184.050 132.760 199.330 ;
        RECT 133.240 196.690 133.590 198.850 ;
        RECT 133.240 184.530 133.590 186.690 ;
        RECT 134.070 184.050 134.240 199.330 ;
        RECT 142.500 198.720 144.480 199.410 ;
        RECT 132.590 183.880 134.240 184.050 ;
        RECT 136.340 198.550 144.480 198.720 ;
        RECT 136.340 184.140 136.510 198.550 ;
        RECT 137.235 197.980 141.775 198.150 ;
        RECT 136.850 197.570 137.020 197.920 ;
        RECT 141.990 197.570 142.160 197.920 ;
        RECT 142.500 197.560 144.480 198.550 ;
        RECT 144.815 198.115 144.995 198.935 ;
        RECT 145.205 198.920 146.745 199.090 ;
        RECT 145.205 198.440 146.745 198.610 ;
        RECT 145.205 197.960 146.745 198.130 ;
        RECT 146.955 198.115 147.135 198.935 ;
        RECT 147.470 197.560 147.640 199.490 ;
        RECT 151.260 199.140 152.920 199.410 ;
        RECT 137.235 197.340 141.775 197.510 ;
        RECT 142.500 197.390 147.640 197.560 ;
        RECT 136.850 196.930 137.020 197.280 ;
        RECT 141.990 196.930 142.160 197.280 ;
        RECT 137.235 196.700 141.775 196.870 ;
        RECT 136.850 196.290 137.020 196.640 ;
        RECT 141.990 196.290 142.160 196.640 ;
        RECT 137.235 196.060 141.775 196.230 ;
        RECT 136.850 195.650 137.020 196.000 ;
        RECT 141.990 195.650 142.160 196.000 ;
        RECT 137.235 195.420 141.775 195.590 ;
        RECT 142.500 195.460 144.480 197.390 ;
        RECT 144.815 196.015 144.995 196.835 ;
        RECT 145.205 196.820 146.745 196.990 ;
        RECT 145.205 196.340 146.745 196.510 ;
        RECT 145.205 195.860 146.745 196.030 ;
        RECT 146.955 196.015 147.135 196.835 ;
        RECT 147.470 195.460 147.640 197.390 ;
        RECT 148.200 198.970 152.920 199.140 ;
        RECT 148.200 197.560 148.370 198.970 ;
        RECT 148.710 198.100 148.880 198.430 ;
        RECT 149.050 198.400 150.590 198.570 ;
        RECT 149.050 197.960 150.590 198.130 ;
        RECT 150.760 198.100 150.930 198.430 ;
        RECT 151.260 197.560 152.920 198.970 ;
        RECT 148.200 197.390 152.920 197.560 ;
        RECT 148.200 195.980 148.370 197.390 ;
        RECT 148.710 196.520 148.880 196.850 ;
        RECT 149.050 196.820 150.590 196.990 ;
        RECT 149.050 196.380 150.590 196.550 ;
        RECT 150.760 196.520 150.930 196.850 ;
        RECT 151.260 195.980 152.920 197.390 ;
        RECT 148.200 195.810 152.920 195.980 ;
        RECT 136.850 195.010 137.020 195.360 ;
        RECT 141.990 195.010 142.160 195.360 ;
        RECT 142.500 195.290 147.640 195.460 ;
        RECT 137.235 194.780 141.775 194.950 ;
        RECT 136.850 194.370 137.020 194.720 ;
        RECT 141.990 194.370 142.160 194.720 ;
        RECT 137.235 194.140 141.775 194.310 ;
        RECT 136.850 193.730 137.020 194.080 ;
        RECT 141.990 193.730 142.160 194.080 ;
        RECT 137.235 193.500 141.775 193.670 ;
        RECT 136.850 193.090 137.020 193.440 ;
        RECT 141.990 193.090 142.160 193.440 ;
        RECT 137.235 192.860 141.775 193.030 ;
        RECT 136.850 192.450 137.020 192.800 ;
        RECT 141.990 192.450 142.160 192.800 ;
        RECT 137.235 192.220 141.775 192.390 ;
        RECT 136.850 191.810 137.020 192.160 ;
        RECT 141.990 191.810 142.160 192.160 ;
        RECT 137.235 191.580 141.775 191.750 ;
        RECT 136.850 191.170 137.020 191.520 ;
        RECT 141.990 191.170 142.160 191.520 ;
        RECT 137.235 190.940 141.775 191.110 ;
        RECT 136.850 190.530 137.020 190.880 ;
        RECT 141.990 190.530 142.160 190.880 ;
        RECT 137.235 190.300 141.775 190.470 ;
        RECT 136.850 189.890 137.020 190.240 ;
        RECT 141.990 189.890 142.160 190.240 ;
        RECT 137.235 189.660 141.775 189.830 ;
        RECT 136.850 189.250 137.020 189.600 ;
        RECT 141.990 189.250 142.160 189.600 ;
        RECT 137.235 189.020 141.775 189.190 ;
        RECT 136.850 188.610 137.020 188.960 ;
        RECT 141.990 188.610 142.160 188.960 ;
        RECT 137.235 188.380 141.775 188.550 ;
        RECT 136.850 187.970 137.020 188.320 ;
        RECT 141.990 187.970 142.160 188.320 ;
        RECT 137.235 187.740 141.775 187.910 ;
        RECT 136.850 187.330 137.020 187.680 ;
        RECT 141.990 187.330 142.160 187.680 ;
        RECT 137.235 187.100 141.775 187.270 ;
        RECT 136.850 186.690 137.020 187.040 ;
        RECT 141.990 186.690 142.160 187.040 ;
        RECT 137.235 186.460 141.775 186.630 ;
        RECT 136.850 186.050 137.020 186.400 ;
        RECT 141.990 186.050 142.160 186.400 ;
        RECT 137.235 185.820 141.775 185.990 ;
        RECT 136.850 185.410 137.020 185.760 ;
        RECT 141.990 185.410 142.160 185.760 ;
        RECT 137.235 185.180 141.775 185.350 ;
        RECT 136.850 184.770 137.020 185.120 ;
        RECT 141.990 184.770 142.160 185.120 ;
        RECT 137.235 184.540 141.775 184.710 ;
        RECT 142.500 184.140 144.120 195.290 ;
        RECT 151.260 193.700 152.920 195.810 ;
        RECT 144.800 193.530 152.920 193.700 ;
        RECT 144.800 188.080 144.970 193.530 ;
        RECT 145.650 192.960 150.190 193.130 ;
        RECT 145.310 192.550 145.480 192.900 ;
        RECT 150.360 192.550 150.530 192.900 ;
        RECT 145.650 192.320 150.190 192.490 ;
        RECT 145.310 191.910 145.480 192.260 ;
        RECT 150.360 191.910 150.530 192.260 ;
        RECT 145.650 191.680 150.190 191.850 ;
        RECT 145.310 191.270 145.480 191.620 ;
        RECT 150.360 191.270 150.530 191.620 ;
        RECT 145.650 191.040 150.190 191.210 ;
        RECT 145.310 190.630 145.480 190.980 ;
        RECT 150.360 190.630 150.530 190.980 ;
        RECT 145.650 190.400 150.190 190.570 ;
        RECT 145.310 189.990 145.480 190.340 ;
        RECT 150.360 189.990 150.530 190.340 ;
        RECT 145.650 189.760 150.190 189.930 ;
        RECT 145.310 189.350 145.480 189.700 ;
        RECT 150.360 189.350 150.530 189.700 ;
        RECT 145.650 189.120 150.190 189.290 ;
        RECT 145.310 188.710 145.480 189.060 ;
        RECT 150.360 188.710 150.530 189.060 ;
        RECT 145.650 188.480 150.190 188.650 ;
        RECT 150.870 188.080 152.920 193.530 ;
        RECT 144.800 187.910 152.920 188.080 ;
        RECT 136.340 183.970 144.120 184.140 ;
        RECT 142.500 182.210 144.120 183.970 ;
        RECT 151.720 182.210 152.920 187.910 ;
        RECT 61.340 173.510 62.030 173.520 ;
        RECT 60.860 173.340 62.510 173.510 ;
        RECT 72.580 173.500 75.910 173.670 ;
        RECT 107.420 173.620 108.110 173.630 ;
        RECT 72.580 173.420 72.750 173.500 ;
        RECT 60.860 158.060 61.030 173.340 ;
        RECT 61.510 170.700 61.860 172.860 ;
        RECT 61.510 158.540 61.860 160.700 ;
        RECT 62.340 158.060 62.510 173.340 ;
        RECT 70.770 172.730 72.750 173.420 ;
        RECT 60.860 157.890 62.510 158.060 ;
        RECT 64.610 172.560 72.750 172.730 ;
        RECT 64.610 158.150 64.780 172.560 ;
        RECT 65.505 171.990 70.045 172.160 ;
        RECT 65.120 171.580 65.290 171.930 ;
        RECT 70.260 171.580 70.430 171.930 ;
        RECT 70.770 171.570 72.750 172.560 ;
        RECT 73.085 172.125 73.265 172.945 ;
        RECT 73.475 172.930 75.015 173.100 ;
        RECT 73.475 172.450 75.015 172.620 ;
        RECT 73.475 171.970 75.015 172.140 ;
        RECT 75.225 172.125 75.405 172.945 ;
        RECT 75.740 171.570 75.910 173.500 ;
        RECT 84.520 173.420 85.210 173.430 ;
        RECT 79.530 173.150 81.190 173.420 ;
        RECT 65.505 171.350 70.045 171.520 ;
        RECT 70.770 171.400 75.910 171.570 ;
        RECT 65.120 170.940 65.290 171.290 ;
        RECT 70.260 170.940 70.430 171.290 ;
        RECT 65.505 170.710 70.045 170.880 ;
        RECT 65.120 170.300 65.290 170.650 ;
        RECT 70.260 170.300 70.430 170.650 ;
        RECT 65.505 170.070 70.045 170.240 ;
        RECT 65.120 169.660 65.290 170.010 ;
        RECT 70.260 169.660 70.430 170.010 ;
        RECT 65.505 169.430 70.045 169.600 ;
        RECT 70.770 169.470 72.750 171.400 ;
        RECT 73.085 170.025 73.265 170.845 ;
        RECT 73.475 170.830 75.015 171.000 ;
        RECT 73.475 170.350 75.015 170.520 ;
        RECT 73.475 169.870 75.015 170.040 ;
        RECT 75.225 170.025 75.405 170.845 ;
        RECT 75.740 169.470 75.910 171.400 ;
        RECT 76.470 172.980 81.190 173.150 ;
        RECT 76.470 171.570 76.640 172.980 ;
        RECT 76.980 172.110 77.150 172.440 ;
        RECT 77.320 172.410 78.860 172.580 ;
        RECT 77.320 171.970 78.860 172.140 ;
        RECT 79.030 172.110 79.200 172.440 ;
        RECT 79.530 171.570 81.190 172.980 ;
        RECT 76.470 171.400 81.190 171.570 ;
        RECT 76.470 169.990 76.640 171.400 ;
        RECT 76.980 170.530 77.150 170.860 ;
        RECT 77.320 170.830 78.860 171.000 ;
        RECT 77.320 170.390 78.860 170.560 ;
        RECT 79.030 170.530 79.200 170.860 ;
        RECT 79.530 169.990 81.190 171.400 ;
        RECT 76.470 169.820 81.190 169.990 ;
        RECT 65.120 169.020 65.290 169.370 ;
        RECT 70.260 169.020 70.430 169.370 ;
        RECT 70.770 169.300 75.910 169.470 ;
        RECT 65.505 168.790 70.045 168.960 ;
        RECT 65.120 168.380 65.290 168.730 ;
        RECT 70.260 168.380 70.430 168.730 ;
        RECT 65.505 168.150 70.045 168.320 ;
        RECT 65.120 167.740 65.290 168.090 ;
        RECT 70.260 167.740 70.430 168.090 ;
        RECT 65.505 167.510 70.045 167.680 ;
        RECT 65.120 167.100 65.290 167.450 ;
        RECT 70.260 167.100 70.430 167.450 ;
        RECT 65.505 166.870 70.045 167.040 ;
        RECT 65.120 166.460 65.290 166.810 ;
        RECT 70.260 166.460 70.430 166.810 ;
        RECT 65.505 166.230 70.045 166.400 ;
        RECT 65.120 165.820 65.290 166.170 ;
        RECT 70.260 165.820 70.430 166.170 ;
        RECT 65.505 165.590 70.045 165.760 ;
        RECT 65.120 165.180 65.290 165.530 ;
        RECT 70.260 165.180 70.430 165.530 ;
        RECT 65.505 164.950 70.045 165.120 ;
        RECT 65.120 164.540 65.290 164.890 ;
        RECT 70.260 164.540 70.430 164.890 ;
        RECT 65.505 164.310 70.045 164.480 ;
        RECT 65.120 163.900 65.290 164.250 ;
        RECT 70.260 163.900 70.430 164.250 ;
        RECT 65.505 163.670 70.045 163.840 ;
        RECT 65.120 163.260 65.290 163.610 ;
        RECT 70.260 163.260 70.430 163.610 ;
        RECT 65.505 163.030 70.045 163.200 ;
        RECT 65.120 162.620 65.290 162.970 ;
        RECT 70.260 162.620 70.430 162.970 ;
        RECT 65.505 162.390 70.045 162.560 ;
        RECT 65.120 161.980 65.290 162.330 ;
        RECT 70.260 161.980 70.430 162.330 ;
        RECT 65.505 161.750 70.045 161.920 ;
        RECT 65.120 161.340 65.290 161.690 ;
        RECT 70.260 161.340 70.430 161.690 ;
        RECT 65.505 161.110 70.045 161.280 ;
        RECT 65.120 160.700 65.290 161.050 ;
        RECT 70.260 160.700 70.430 161.050 ;
        RECT 65.505 160.470 70.045 160.640 ;
        RECT 65.120 160.060 65.290 160.410 ;
        RECT 70.260 160.060 70.430 160.410 ;
        RECT 65.505 159.830 70.045 160.000 ;
        RECT 65.120 159.420 65.290 159.770 ;
        RECT 70.260 159.420 70.430 159.770 ;
        RECT 65.505 159.190 70.045 159.360 ;
        RECT 65.120 158.780 65.290 159.130 ;
        RECT 70.260 158.780 70.430 159.130 ;
        RECT 65.505 158.550 70.045 158.720 ;
        RECT 70.770 158.150 72.390 169.300 ;
        RECT 79.530 167.710 81.190 169.820 ;
        RECT 73.070 167.540 81.190 167.710 ;
        RECT 73.070 162.090 73.240 167.540 ;
        RECT 73.920 166.970 78.460 167.140 ;
        RECT 73.580 166.560 73.750 166.910 ;
        RECT 78.630 166.560 78.800 166.910 ;
        RECT 73.920 166.330 78.460 166.500 ;
        RECT 73.580 165.920 73.750 166.270 ;
        RECT 78.630 165.920 78.800 166.270 ;
        RECT 73.920 165.690 78.460 165.860 ;
        RECT 73.580 165.280 73.750 165.630 ;
        RECT 78.630 165.280 78.800 165.630 ;
        RECT 73.920 165.050 78.460 165.220 ;
        RECT 73.580 164.640 73.750 164.990 ;
        RECT 78.630 164.640 78.800 164.990 ;
        RECT 73.920 164.410 78.460 164.580 ;
        RECT 73.580 164.000 73.750 164.350 ;
        RECT 78.630 164.000 78.800 164.350 ;
        RECT 73.920 163.770 78.460 163.940 ;
        RECT 73.580 163.360 73.750 163.710 ;
        RECT 78.630 163.360 78.800 163.710 ;
        RECT 73.920 163.130 78.460 163.300 ;
        RECT 73.580 162.720 73.750 163.070 ;
        RECT 78.630 162.720 78.800 163.070 ;
        RECT 73.920 162.490 78.460 162.660 ;
        RECT 79.140 162.090 81.190 167.540 ;
        RECT 73.070 161.920 81.190 162.090 ;
        RECT 64.610 157.980 72.390 158.150 ;
        RECT 70.770 156.220 72.390 157.980 ;
        RECT 79.990 156.220 81.190 161.920 ;
        RECT 84.040 173.250 85.690 173.420 ;
        RECT 95.760 173.410 99.090 173.580 ;
        RECT 95.760 173.330 95.930 173.410 ;
        RECT 84.040 157.970 84.210 173.250 ;
        RECT 84.690 170.610 85.040 172.770 ;
        RECT 84.690 158.450 85.040 160.610 ;
        RECT 85.520 157.970 85.690 173.250 ;
        RECT 93.950 172.640 95.930 173.330 ;
        RECT 84.040 157.800 85.690 157.970 ;
        RECT 87.790 172.470 95.930 172.640 ;
        RECT 87.790 158.060 87.960 172.470 ;
        RECT 88.685 171.900 93.225 172.070 ;
        RECT 88.300 171.490 88.470 171.840 ;
        RECT 93.440 171.490 93.610 171.840 ;
        RECT 93.950 171.480 95.930 172.470 ;
        RECT 96.265 172.035 96.445 172.855 ;
        RECT 96.655 172.840 98.195 173.010 ;
        RECT 96.655 172.360 98.195 172.530 ;
        RECT 96.655 171.880 98.195 172.050 ;
        RECT 98.405 172.035 98.585 172.855 ;
        RECT 98.920 171.480 99.090 173.410 ;
        RECT 106.940 173.450 108.590 173.620 ;
        RECT 118.660 173.610 121.990 173.780 ;
        RECT 130.520 173.730 131.210 173.740 ;
        RECT 118.660 173.530 118.830 173.610 ;
        RECT 102.710 173.060 104.370 173.330 ;
        RECT 88.685 171.260 93.225 171.430 ;
        RECT 93.950 171.310 99.090 171.480 ;
        RECT 88.300 170.850 88.470 171.200 ;
        RECT 93.440 170.850 93.610 171.200 ;
        RECT 88.685 170.620 93.225 170.790 ;
        RECT 88.300 170.210 88.470 170.560 ;
        RECT 93.440 170.210 93.610 170.560 ;
        RECT 88.685 169.980 93.225 170.150 ;
        RECT 88.300 169.570 88.470 169.920 ;
        RECT 93.440 169.570 93.610 169.920 ;
        RECT 88.685 169.340 93.225 169.510 ;
        RECT 93.950 169.380 95.930 171.310 ;
        RECT 96.265 169.935 96.445 170.755 ;
        RECT 96.655 170.740 98.195 170.910 ;
        RECT 96.655 170.260 98.195 170.430 ;
        RECT 96.655 169.780 98.195 169.950 ;
        RECT 98.405 169.935 98.585 170.755 ;
        RECT 98.920 169.380 99.090 171.310 ;
        RECT 99.650 172.890 104.370 173.060 ;
        RECT 99.650 171.480 99.820 172.890 ;
        RECT 100.160 172.020 100.330 172.350 ;
        RECT 100.500 172.320 102.040 172.490 ;
        RECT 100.500 171.880 102.040 172.050 ;
        RECT 102.210 172.020 102.380 172.350 ;
        RECT 102.710 171.480 104.370 172.890 ;
        RECT 99.650 171.310 104.370 171.480 ;
        RECT 99.650 169.900 99.820 171.310 ;
        RECT 100.160 170.440 100.330 170.770 ;
        RECT 100.500 170.740 102.040 170.910 ;
        RECT 100.500 170.300 102.040 170.470 ;
        RECT 102.210 170.440 102.380 170.770 ;
        RECT 102.710 169.900 104.370 171.310 ;
        RECT 99.650 169.730 104.370 169.900 ;
        RECT 88.300 168.930 88.470 169.280 ;
        RECT 93.440 168.930 93.610 169.280 ;
        RECT 93.950 169.210 99.090 169.380 ;
        RECT 88.685 168.700 93.225 168.870 ;
        RECT 88.300 168.290 88.470 168.640 ;
        RECT 93.440 168.290 93.610 168.640 ;
        RECT 88.685 168.060 93.225 168.230 ;
        RECT 88.300 167.650 88.470 168.000 ;
        RECT 93.440 167.650 93.610 168.000 ;
        RECT 88.685 167.420 93.225 167.590 ;
        RECT 88.300 167.010 88.470 167.360 ;
        RECT 93.440 167.010 93.610 167.360 ;
        RECT 88.685 166.780 93.225 166.950 ;
        RECT 88.300 166.370 88.470 166.720 ;
        RECT 93.440 166.370 93.610 166.720 ;
        RECT 88.685 166.140 93.225 166.310 ;
        RECT 88.300 165.730 88.470 166.080 ;
        RECT 93.440 165.730 93.610 166.080 ;
        RECT 88.685 165.500 93.225 165.670 ;
        RECT 88.300 165.090 88.470 165.440 ;
        RECT 93.440 165.090 93.610 165.440 ;
        RECT 88.685 164.860 93.225 165.030 ;
        RECT 88.300 164.450 88.470 164.800 ;
        RECT 93.440 164.450 93.610 164.800 ;
        RECT 88.685 164.220 93.225 164.390 ;
        RECT 88.300 163.810 88.470 164.160 ;
        RECT 93.440 163.810 93.610 164.160 ;
        RECT 88.685 163.580 93.225 163.750 ;
        RECT 88.300 163.170 88.470 163.520 ;
        RECT 93.440 163.170 93.610 163.520 ;
        RECT 88.685 162.940 93.225 163.110 ;
        RECT 88.300 162.530 88.470 162.880 ;
        RECT 93.440 162.530 93.610 162.880 ;
        RECT 88.685 162.300 93.225 162.470 ;
        RECT 88.300 161.890 88.470 162.240 ;
        RECT 93.440 161.890 93.610 162.240 ;
        RECT 88.685 161.660 93.225 161.830 ;
        RECT 88.300 161.250 88.470 161.600 ;
        RECT 93.440 161.250 93.610 161.600 ;
        RECT 88.685 161.020 93.225 161.190 ;
        RECT 88.300 160.610 88.470 160.960 ;
        RECT 93.440 160.610 93.610 160.960 ;
        RECT 88.685 160.380 93.225 160.550 ;
        RECT 88.300 159.970 88.470 160.320 ;
        RECT 93.440 159.970 93.610 160.320 ;
        RECT 88.685 159.740 93.225 159.910 ;
        RECT 88.300 159.330 88.470 159.680 ;
        RECT 93.440 159.330 93.610 159.680 ;
        RECT 88.685 159.100 93.225 159.270 ;
        RECT 88.300 158.690 88.470 159.040 ;
        RECT 93.440 158.690 93.610 159.040 ;
        RECT 88.685 158.460 93.225 158.630 ;
        RECT 93.950 158.060 95.570 169.210 ;
        RECT 102.710 167.620 104.370 169.730 ;
        RECT 96.250 167.450 104.370 167.620 ;
        RECT 96.250 162.000 96.420 167.450 ;
        RECT 97.100 166.880 101.640 167.050 ;
        RECT 96.760 166.470 96.930 166.820 ;
        RECT 101.810 166.470 101.980 166.820 ;
        RECT 97.100 166.240 101.640 166.410 ;
        RECT 96.760 165.830 96.930 166.180 ;
        RECT 101.810 165.830 101.980 166.180 ;
        RECT 97.100 165.600 101.640 165.770 ;
        RECT 96.760 165.190 96.930 165.540 ;
        RECT 101.810 165.190 101.980 165.540 ;
        RECT 97.100 164.960 101.640 165.130 ;
        RECT 96.760 164.550 96.930 164.900 ;
        RECT 101.810 164.550 101.980 164.900 ;
        RECT 97.100 164.320 101.640 164.490 ;
        RECT 96.760 163.910 96.930 164.260 ;
        RECT 101.810 163.910 101.980 164.260 ;
        RECT 97.100 163.680 101.640 163.850 ;
        RECT 96.760 163.270 96.930 163.620 ;
        RECT 101.810 163.270 101.980 163.620 ;
        RECT 97.100 163.040 101.640 163.210 ;
        RECT 96.760 162.630 96.930 162.980 ;
        RECT 101.810 162.630 101.980 162.980 ;
        RECT 97.100 162.400 101.640 162.570 ;
        RECT 102.320 162.000 104.370 167.450 ;
        RECT 96.250 161.830 104.370 162.000 ;
        RECT 87.790 157.890 95.570 158.060 ;
        RECT 93.950 156.130 95.570 157.890 ;
        RECT 103.170 156.130 104.370 161.830 ;
        RECT 106.940 158.170 107.110 173.450 ;
        RECT 107.590 170.810 107.940 172.970 ;
        RECT 107.590 158.650 107.940 160.810 ;
        RECT 108.420 158.170 108.590 173.450 ;
        RECT 116.850 172.840 118.830 173.530 ;
        RECT 106.940 158.000 108.590 158.170 ;
        RECT 110.690 172.670 118.830 172.840 ;
        RECT 110.690 158.260 110.860 172.670 ;
        RECT 111.585 172.100 116.125 172.270 ;
        RECT 111.200 171.690 111.370 172.040 ;
        RECT 116.340 171.690 116.510 172.040 ;
        RECT 116.850 171.680 118.830 172.670 ;
        RECT 119.165 172.235 119.345 173.055 ;
        RECT 119.555 173.040 121.095 173.210 ;
        RECT 119.555 172.560 121.095 172.730 ;
        RECT 119.555 172.080 121.095 172.250 ;
        RECT 121.305 172.235 121.485 173.055 ;
        RECT 121.820 171.680 121.990 173.610 ;
        RECT 130.040 173.560 131.690 173.730 ;
        RECT 141.760 173.720 145.090 173.890 ;
        RECT 141.760 173.640 141.930 173.720 ;
        RECT 125.610 173.260 127.270 173.530 ;
        RECT 111.585 171.460 116.125 171.630 ;
        RECT 116.850 171.510 121.990 171.680 ;
        RECT 111.200 171.050 111.370 171.400 ;
        RECT 116.340 171.050 116.510 171.400 ;
        RECT 111.585 170.820 116.125 170.990 ;
        RECT 111.200 170.410 111.370 170.760 ;
        RECT 116.340 170.410 116.510 170.760 ;
        RECT 111.585 170.180 116.125 170.350 ;
        RECT 111.200 169.770 111.370 170.120 ;
        RECT 116.340 169.770 116.510 170.120 ;
        RECT 111.585 169.540 116.125 169.710 ;
        RECT 116.850 169.580 118.830 171.510 ;
        RECT 119.165 170.135 119.345 170.955 ;
        RECT 119.555 170.940 121.095 171.110 ;
        RECT 119.555 170.460 121.095 170.630 ;
        RECT 119.555 169.980 121.095 170.150 ;
        RECT 121.305 170.135 121.485 170.955 ;
        RECT 121.820 169.580 121.990 171.510 ;
        RECT 122.550 173.090 127.270 173.260 ;
        RECT 122.550 171.680 122.720 173.090 ;
        RECT 123.060 172.220 123.230 172.550 ;
        RECT 123.400 172.520 124.940 172.690 ;
        RECT 123.400 172.080 124.940 172.250 ;
        RECT 125.110 172.220 125.280 172.550 ;
        RECT 125.610 171.680 127.270 173.090 ;
        RECT 122.550 171.510 127.270 171.680 ;
        RECT 122.550 170.100 122.720 171.510 ;
        RECT 123.060 170.640 123.230 170.970 ;
        RECT 123.400 170.940 124.940 171.110 ;
        RECT 123.400 170.500 124.940 170.670 ;
        RECT 125.110 170.640 125.280 170.970 ;
        RECT 125.610 170.100 127.270 171.510 ;
        RECT 122.550 169.930 127.270 170.100 ;
        RECT 111.200 169.130 111.370 169.480 ;
        RECT 116.340 169.130 116.510 169.480 ;
        RECT 116.850 169.410 121.990 169.580 ;
        RECT 111.585 168.900 116.125 169.070 ;
        RECT 111.200 168.490 111.370 168.840 ;
        RECT 116.340 168.490 116.510 168.840 ;
        RECT 111.585 168.260 116.125 168.430 ;
        RECT 111.200 167.850 111.370 168.200 ;
        RECT 116.340 167.850 116.510 168.200 ;
        RECT 111.585 167.620 116.125 167.790 ;
        RECT 111.200 167.210 111.370 167.560 ;
        RECT 116.340 167.210 116.510 167.560 ;
        RECT 111.585 166.980 116.125 167.150 ;
        RECT 111.200 166.570 111.370 166.920 ;
        RECT 116.340 166.570 116.510 166.920 ;
        RECT 111.585 166.340 116.125 166.510 ;
        RECT 111.200 165.930 111.370 166.280 ;
        RECT 116.340 165.930 116.510 166.280 ;
        RECT 111.585 165.700 116.125 165.870 ;
        RECT 111.200 165.290 111.370 165.640 ;
        RECT 116.340 165.290 116.510 165.640 ;
        RECT 111.585 165.060 116.125 165.230 ;
        RECT 111.200 164.650 111.370 165.000 ;
        RECT 116.340 164.650 116.510 165.000 ;
        RECT 111.585 164.420 116.125 164.590 ;
        RECT 111.200 164.010 111.370 164.360 ;
        RECT 116.340 164.010 116.510 164.360 ;
        RECT 111.585 163.780 116.125 163.950 ;
        RECT 111.200 163.370 111.370 163.720 ;
        RECT 116.340 163.370 116.510 163.720 ;
        RECT 111.585 163.140 116.125 163.310 ;
        RECT 111.200 162.730 111.370 163.080 ;
        RECT 116.340 162.730 116.510 163.080 ;
        RECT 111.585 162.500 116.125 162.670 ;
        RECT 111.200 162.090 111.370 162.440 ;
        RECT 116.340 162.090 116.510 162.440 ;
        RECT 111.585 161.860 116.125 162.030 ;
        RECT 111.200 161.450 111.370 161.800 ;
        RECT 116.340 161.450 116.510 161.800 ;
        RECT 111.585 161.220 116.125 161.390 ;
        RECT 111.200 160.810 111.370 161.160 ;
        RECT 116.340 160.810 116.510 161.160 ;
        RECT 111.585 160.580 116.125 160.750 ;
        RECT 111.200 160.170 111.370 160.520 ;
        RECT 116.340 160.170 116.510 160.520 ;
        RECT 111.585 159.940 116.125 160.110 ;
        RECT 111.200 159.530 111.370 159.880 ;
        RECT 116.340 159.530 116.510 159.880 ;
        RECT 111.585 159.300 116.125 159.470 ;
        RECT 111.200 158.890 111.370 159.240 ;
        RECT 116.340 158.890 116.510 159.240 ;
        RECT 111.585 158.660 116.125 158.830 ;
        RECT 116.850 158.260 118.470 169.410 ;
        RECT 125.610 167.820 127.270 169.930 ;
        RECT 119.150 167.650 127.270 167.820 ;
        RECT 119.150 162.200 119.320 167.650 ;
        RECT 120.000 167.080 124.540 167.250 ;
        RECT 119.660 166.670 119.830 167.020 ;
        RECT 124.710 166.670 124.880 167.020 ;
        RECT 120.000 166.440 124.540 166.610 ;
        RECT 119.660 166.030 119.830 166.380 ;
        RECT 124.710 166.030 124.880 166.380 ;
        RECT 120.000 165.800 124.540 165.970 ;
        RECT 119.660 165.390 119.830 165.740 ;
        RECT 124.710 165.390 124.880 165.740 ;
        RECT 120.000 165.160 124.540 165.330 ;
        RECT 119.660 164.750 119.830 165.100 ;
        RECT 124.710 164.750 124.880 165.100 ;
        RECT 120.000 164.520 124.540 164.690 ;
        RECT 119.660 164.110 119.830 164.460 ;
        RECT 124.710 164.110 124.880 164.460 ;
        RECT 120.000 163.880 124.540 164.050 ;
        RECT 119.660 163.470 119.830 163.820 ;
        RECT 124.710 163.470 124.880 163.820 ;
        RECT 120.000 163.240 124.540 163.410 ;
        RECT 119.660 162.830 119.830 163.180 ;
        RECT 124.710 162.830 124.880 163.180 ;
        RECT 120.000 162.600 124.540 162.770 ;
        RECT 125.220 162.200 127.270 167.650 ;
        RECT 119.150 162.030 127.270 162.200 ;
        RECT 110.690 158.090 118.470 158.260 ;
        RECT 116.850 156.330 118.470 158.090 ;
        RECT 126.070 156.330 127.270 162.030 ;
        RECT 130.040 158.280 130.210 173.560 ;
        RECT 130.690 170.920 131.040 173.080 ;
        RECT 130.690 158.760 131.040 160.920 ;
        RECT 131.520 158.280 131.690 173.560 ;
        RECT 139.950 172.950 141.930 173.640 ;
        RECT 130.040 158.110 131.690 158.280 ;
        RECT 133.790 172.780 141.930 172.950 ;
        RECT 133.790 158.370 133.960 172.780 ;
        RECT 134.685 172.210 139.225 172.380 ;
        RECT 134.300 171.800 134.470 172.150 ;
        RECT 139.440 171.800 139.610 172.150 ;
        RECT 139.950 171.790 141.930 172.780 ;
        RECT 142.265 172.345 142.445 173.165 ;
        RECT 142.655 173.150 144.195 173.320 ;
        RECT 142.655 172.670 144.195 172.840 ;
        RECT 142.655 172.190 144.195 172.360 ;
        RECT 144.405 172.345 144.585 173.165 ;
        RECT 144.920 171.790 145.090 173.720 ;
        RECT 148.710 173.370 150.370 173.640 ;
        RECT 134.685 171.570 139.225 171.740 ;
        RECT 139.950 171.620 145.090 171.790 ;
        RECT 134.300 171.160 134.470 171.510 ;
        RECT 139.440 171.160 139.610 171.510 ;
        RECT 134.685 170.930 139.225 171.100 ;
        RECT 134.300 170.520 134.470 170.870 ;
        RECT 139.440 170.520 139.610 170.870 ;
        RECT 134.685 170.290 139.225 170.460 ;
        RECT 134.300 169.880 134.470 170.230 ;
        RECT 139.440 169.880 139.610 170.230 ;
        RECT 134.685 169.650 139.225 169.820 ;
        RECT 139.950 169.690 141.930 171.620 ;
        RECT 142.265 170.245 142.445 171.065 ;
        RECT 142.655 171.050 144.195 171.220 ;
        RECT 142.655 170.570 144.195 170.740 ;
        RECT 142.655 170.090 144.195 170.260 ;
        RECT 144.405 170.245 144.585 171.065 ;
        RECT 144.920 169.690 145.090 171.620 ;
        RECT 145.650 173.200 150.370 173.370 ;
        RECT 145.650 171.790 145.820 173.200 ;
        RECT 146.160 172.330 146.330 172.660 ;
        RECT 146.500 172.630 148.040 172.800 ;
        RECT 146.500 172.190 148.040 172.360 ;
        RECT 148.210 172.330 148.380 172.660 ;
        RECT 148.710 171.790 150.370 173.200 ;
        RECT 145.650 171.620 150.370 171.790 ;
        RECT 145.650 170.210 145.820 171.620 ;
        RECT 146.160 170.750 146.330 171.080 ;
        RECT 146.500 171.050 148.040 171.220 ;
        RECT 146.500 170.610 148.040 170.780 ;
        RECT 148.210 170.750 148.380 171.080 ;
        RECT 148.710 170.210 150.370 171.620 ;
        RECT 145.650 170.040 150.370 170.210 ;
        RECT 134.300 169.240 134.470 169.590 ;
        RECT 139.440 169.240 139.610 169.590 ;
        RECT 139.950 169.520 145.090 169.690 ;
        RECT 134.685 169.010 139.225 169.180 ;
        RECT 134.300 168.600 134.470 168.950 ;
        RECT 139.440 168.600 139.610 168.950 ;
        RECT 134.685 168.370 139.225 168.540 ;
        RECT 134.300 167.960 134.470 168.310 ;
        RECT 139.440 167.960 139.610 168.310 ;
        RECT 134.685 167.730 139.225 167.900 ;
        RECT 134.300 167.320 134.470 167.670 ;
        RECT 139.440 167.320 139.610 167.670 ;
        RECT 134.685 167.090 139.225 167.260 ;
        RECT 134.300 166.680 134.470 167.030 ;
        RECT 139.440 166.680 139.610 167.030 ;
        RECT 134.685 166.450 139.225 166.620 ;
        RECT 134.300 166.040 134.470 166.390 ;
        RECT 139.440 166.040 139.610 166.390 ;
        RECT 134.685 165.810 139.225 165.980 ;
        RECT 134.300 165.400 134.470 165.750 ;
        RECT 139.440 165.400 139.610 165.750 ;
        RECT 134.685 165.170 139.225 165.340 ;
        RECT 134.300 164.760 134.470 165.110 ;
        RECT 139.440 164.760 139.610 165.110 ;
        RECT 134.685 164.530 139.225 164.700 ;
        RECT 134.300 164.120 134.470 164.470 ;
        RECT 139.440 164.120 139.610 164.470 ;
        RECT 134.685 163.890 139.225 164.060 ;
        RECT 134.300 163.480 134.470 163.830 ;
        RECT 139.440 163.480 139.610 163.830 ;
        RECT 134.685 163.250 139.225 163.420 ;
        RECT 134.300 162.840 134.470 163.190 ;
        RECT 139.440 162.840 139.610 163.190 ;
        RECT 134.685 162.610 139.225 162.780 ;
        RECT 134.300 162.200 134.470 162.550 ;
        RECT 139.440 162.200 139.610 162.550 ;
        RECT 134.685 161.970 139.225 162.140 ;
        RECT 134.300 161.560 134.470 161.910 ;
        RECT 139.440 161.560 139.610 161.910 ;
        RECT 134.685 161.330 139.225 161.500 ;
        RECT 134.300 160.920 134.470 161.270 ;
        RECT 139.440 160.920 139.610 161.270 ;
        RECT 134.685 160.690 139.225 160.860 ;
        RECT 134.300 160.280 134.470 160.630 ;
        RECT 139.440 160.280 139.610 160.630 ;
        RECT 134.685 160.050 139.225 160.220 ;
        RECT 134.300 159.640 134.470 159.990 ;
        RECT 139.440 159.640 139.610 159.990 ;
        RECT 134.685 159.410 139.225 159.580 ;
        RECT 134.300 159.000 134.470 159.350 ;
        RECT 139.440 159.000 139.610 159.350 ;
        RECT 134.685 158.770 139.225 158.940 ;
        RECT 139.950 158.370 141.570 169.520 ;
        RECT 148.710 167.930 150.370 170.040 ;
        RECT 142.250 167.760 150.370 167.930 ;
        RECT 142.250 162.310 142.420 167.760 ;
        RECT 143.100 167.190 147.640 167.360 ;
        RECT 142.760 166.780 142.930 167.130 ;
        RECT 147.810 166.780 147.980 167.130 ;
        RECT 143.100 166.550 147.640 166.720 ;
        RECT 142.760 166.140 142.930 166.490 ;
        RECT 147.810 166.140 147.980 166.490 ;
        RECT 143.100 165.910 147.640 166.080 ;
        RECT 142.760 165.500 142.930 165.850 ;
        RECT 147.810 165.500 147.980 165.850 ;
        RECT 143.100 165.270 147.640 165.440 ;
        RECT 142.760 164.860 142.930 165.210 ;
        RECT 147.810 164.860 147.980 165.210 ;
        RECT 143.100 164.630 147.640 164.800 ;
        RECT 142.760 164.220 142.930 164.570 ;
        RECT 147.810 164.220 147.980 164.570 ;
        RECT 143.100 163.990 147.640 164.160 ;
        RECT 142.760 163.580 142.930 163.930 ;
        RECT 147.810 163.580 147.980 163.930 ;
        RECT 143.100 163.350 147.640 163.520 ;
        RECT 142.760 162.940 142.930 163.290 ;
        RECT 147.810 162.940 147.980 163.290 ;
        RECT 143.100 162.710 147.640 162.880 ;
        RECT 148.320 162.310 150.370 167.760 ;
        RECT 142.250 162.140 150.370 162.310 ;
        RECT 133.790 158.200 141.570 158.370 ;
        RECT 139.950 156.440 141.570 158.200 ;
        RECT 149.170 156.440 150.370 162.140 ;
        RECT 84.730 147.780 85.420 147.790 ;
        RECT 84.250 147.610 85.900 147.780 ;
        RECT 95.970 147.770 99.300 147.940 ;
        RECT 107.760 147.930 108.450 147.940 ;
        RECT 95.970 147.690 96.140 147.770 ;
        RECT 84.250 132.330 84.420 147.610 ;
        RECT 84.900 144.970 85.250 147.130 ;
        RECT 84.900 132.810 85.250 134.970 ;
        RECT 85.730 132.330 85.900 147.610 ;
        RECT 94.160 147.000 96.140 147.690 ;
        RECT 84.250 132.160 85.900 132.330 ;
        RECT 88.000 146.830 96.140 147.000 ;
        RECT 88.000 132.420 88.170 146.830 ;
        RECT 88.895 146.260 93.435 146.430 ;
        RECT 88.510 145.850 88.680 146.200 ;
        RECT 93.650 145.850 93.820 146.200 ;
        RECT 94.160 145.840 96.140 146.830 ;
        RECT 96.475 146.395 96.655 147.215 ;
        RECT 96.865 147.200 98.405 147.370 ;
        RECT 96.865 146.720 98.405 146.890 ;
        RECT 96.865 146.240 98.405 146.410 ;
        RECT 98.615 146.395 98.795 147.215 ;
        RECT 99.130 145.840 99.300 147.770 ;
        RECT 107.280 147.760 108.930 147.930 ;
        RECT 119.000 147.920 122.330 148.090 ;
        RECT 130.770 148.010 131.460 148.020 ;
        RECT 119.000 147.840 119.170 147.920 ;
        RECT 102.920 147.420 104.580 147.690 ;
        RECT 88.895 145.620 93.435 145.790 ;
        RECT 94.160 145.670 99.300 145.840 ;
        RECT 88.510 145.210 88.680 145.560 ;
        RECT 93.650 145.210 93.820 145.560 ;
        RECT 88.895 144.980 93.435 145.150 ;
        RECT 88.510 144.570 88.680 144.920 ;
        RECT 93.650 144.570 93.820 144.920 ;
        RECT 88.895 144.340 93.435 144.510 ;
        RECT 88.510 143.930 88.680 144.280 ;
        RECT 93.650 143.930 93.820 144.280 ;
        RECT 88.895 143.700 93.435 143.870 ;
        RECT 94.160 143.740 96.140 145.670 ;
        RECT 96.475 144.295 96.655 145.115 ;
        RECT 96.865 145.100 98.405 145.270 ;
        RECT 96.865 144.620 98.405 144.790 ;
        RECT 96.865 144.140 98.405 144.310 ;
        RECT 98.615 144.295 98.795 145.115 ;
        RECT 99.130 143.740 99.300 145.670 ;
        RECT 99.860 147.250 104.580 147.420 ;
        RECT 99.860 145.840 100.030 147.250 ;
        RECT 100.370 146.380 100.540 146.710 ;
        RECT 100.710 146.680 102.250 146.850 ;
        RECT 100.710 146.240 102.250 146.410 ;
        RECT 102.420 146.380 102.590 146.710 ;
        RECT 102.920 145.840 104.580 147.250 ;
        RECT 99.860 145.670 104.580 145.840 ;
        RECT 99.860 144.260 100.030 145.670 ;
        RECT 100.370 144.800 100.540 145.130 ;
        RECT 100.710 145.100 102.250 145.270 ;
        RECT 100.710 144.660 102.250 144.830 ;
        RECT 102.420 144.800 102.590 145.130 ;
        RECT 102.920 144.260 104.580 145.670 ;
        RECT 99.860 144.090 104.580 144.260 ;
        RECT 88.510 143.290 88.680 143.640 ;
        RECT 93.650 143.290 93.820 143.640 ;
        RECT 94.160 143.570 99.300 143.740 ;
        RECT 88.895 143.060 93.435 143.230 ;
        RECT 88.510 142.650 88.680 143.000 ;
        RECT 93.650 142.650 93.820 143.000 ;
        RECT 88.895 142.420 93.435 142.590 ;
        RECT 88.510 142.010 88.680 142.360 ;
        RECT 93.650 142.010 93.820 142.360 ;
        RECT 88.895 141.780 93.435 141.950 ;
        RECT 88.510 141.370 88.680 141.720 ;
        RECT 93.650 141.370 93.820 141.720 ;
        RECT 88.895 141.140 93.435 141.310 ;
        RECT 88.510 140.730 88.680 141.080 ;
        RECT 93.650 140.730 93.820 141.080 ;
        RECT 88.895 140.500 93.435 140.670 ;
        RECT 88.510 140.090 88.680 140.440 ;
        RECT 93.650 140.090 93.820 140.440 ;
        RECT 88.895 139.860 93.435 140.030 ;
        RECT 88.510 139.450 88.680 139.800 ;
        RECT 93.650 139.450 93.820 139.800 ;
        RECT 88.895 139.220 93.435 139.390 ;
        RECT 88.510 138.810 88.680 139.160 ;
        RECT 93.650 138.810 93.820 139.160 ;
        RECT 88.895 138.580 93.435 138.750 ;
        RECT 88.510 138.170 88.680 138.520 ;
        RECT 93.650 138.170 93.820 138.520 ;
        RECT 88.895 137.940 93.435 138.110 ;
        RECT 88.510 137.530 88.680 137.880 ;
        RECT 93.650 137.530 93.820 137.880 ;
        RECT 88.895 137.300 93.435 137.470 ;
        RECT 88.510 136.890 88.680 137.240 ;
        RECT 93.650 136.890 93.820 137.240 ;
        RECT 88.895 136.660 93.435 136.830 ;
        RECT 88.510 136.250 88.680 136.600 ;
        RECT 93.650 136.250 93.820 136.600 ;
        RECT 88.895 136.020 93.435 136.190 ;
        RECT 88.510 135.610 88.680 135.960 ;
        RECT 93.650 135.610 93.820 135.960 ;
        RECT 88.895 135.380 93.435 135.550 ;
        RECT 88.510 134.970 88.680 135.320 ;
        RECT 93.650 134.970 93.820 135.320 ;
        RECT 88.895 134.740 93.435 134.910 ;
        RECT 88.510 134.330 88.680 134.680 ;
        RECT 93.650 134.330 93.820 134.680 ;
        RECT 88.895 134.100 93.435 134.270 ;
        RECT 88.510 133.690 88.680 134.040 ;
        RECT 93.650 133.690 93.820 134.040 ;
        RECT 88.895 133.460 93.435 133.630 ;
        RECT 88.510 133.050 88.680 133.400 ;
        RECT 93.650 133.050 93.820 133.400 ;
        RECT 88.895 132.820 93.435 132.990 ;
        RECT 94.160 132.420 95.780 143.570 ;
        RECT 102.920 141.980 104.580 144.090 ;
        RECT 96.460 141.810 104.580 141.980 ;
        RECT 96.460 136.360 96.630 141.810 ;
        RECT 97.310 141.240 101.850 141.410 ;
        RECT 96.970 140.830 97.140 141.180 ;
        RECT 102.020 140.830 102.190 141.180 ;
        RECT 97.310 140.600 101.850 140.770 ;
        RECT 96.970 140.190 97.140 140.540 ;
        RECT 102.020 140.190 102.190 140.540 ;
        RECT 97.310 139.960 101.850 140.130 ;
        RECT 96.970 139.550 97.140 139.900 ;
        RECT 102.020 139.550 102.190 139.900 ;
        RECT 97.310 139.320 101.850 139.490 ;
        RECT 96.970 138.910 97.140 139.260 ;
        RECT 102.020 138.910 102.190 139.260 ;
        RECT 97.310 138.680 101.850 138.850 ;
        RECT 96.970 138.270 97.140 138.620 ;
        RECT 102.020 138.270 102.190 138.620 ;
        RECT 97.310 138.040 101.850 138.210 ;
        RECT 96.970 137.630 97.140 137.980 ;
        RECT 102.020 137.630 102.190 137.980 ;
        RECT 97.310 137.400 101.850 137.570 ;
        RECT 96.970 136.990 97.140 137.340 ;
        RECT 102.020 136.990 102.190 137.340 ;
        RECT 97.310 136.760 101.850 136.930 ;
        RECT 102.530 136.360 104.580 141.810 ;
        RECT 96.460 136.190 104.580 136.360 ;
        RECT 88.000 132.250 95.780 132.420 ;
        RECT 94.160 130.490 95.780 132.250 ;
        RECT 103.380 130.490 104.580 136.190 ;
        RECT 107.280 132.480 107.450 147.760 ;
        RECT 107.930 145.120 108.280 147.280 ;
        RECT 107.930 132.960 108.280 135.120 ;
        RECT 108.760 132.480 108.930 147.760 ;
        RECT 117.190 147.150 119.170 147.840 ;
        RECT 107.280 132.310 108.930 132.480 ;
        RECT 111.030 146.980 119.170 147.150 ;
        RECT 111.030 132.570 111.200 146.980 ;
        RECT 111.925 146.410 116.465 146.580 ;
        RECT 111.540 146.000 111.710 146.350 ;
        RECT 116.680 146.000 116.850 146.350 ;
        RECT 117.190 145.990 119.170 146.980 ;
        RECT 119.505 146.545 119.685 147.365 ;
        RECT 119.895 147.350 121.435 147.520 ;
        RECT 119.895 146.870 121.435 147.040 ;
        RECT 119.895 146.390 121.435 146.560 ;
        RECT 121.645 146.545 121.825 147.365 ;
        RECT 122.160 145.990 122.330 147.920 ;
        RECT 130.290 147.840 131.940 148.010 ;
        RECT 142.010 148.000 145.340 148.170 ;
        RECT 142.010 147.920 142.180 148.000 ;
        RECT 125.950 147.570 127.610 147.840 ;
        RECT 111.925 145.770 116.465 145.940 ;
        RECT 117.190 145.820 122.330 145.990 ;
        RECT 111.540 145.360 111.710 145.710 ;
        RECT 116.680 145.360 116.850 145.710 ;
        RECT 111.925 145.130 116.465 145.300 ;
        RECT 111.540 144.720 111.710 145.070 ;
        RECT 116.680 144.720 116.850 145.070 ;
        RECT 111.925 144.490 116.465 144.660 ;
        RECT 111.540 144.080 111.710 144.430 ;
        RECT 116.680 144.080 116.850 144.430 ;
        RECT 111.925 143.850 116.465 144.020 ;
        RECT 117.190 143.890 119.170 145.820 ;
        RECT 119.505 144.445 119.685 145.265 ;
        RECT 119.895 145.250 121.435 145.420 ;
        RECT 119.895 144.770 121.435 144.940 ;
        RECT 119.895 144.290 121.435 144.460 ;
        RECT 121.645 144.445 121.825 145.265 ;
        RECT 122.160 143.890 122.330 145.820 ;
        RECT 122.890 147.400 127.610 147.570 ;
        RECT 122.890 145.990 123.060 147.400 ;
        RECT 123.400 146.530 123.570 146.860 ;
        RECT 123.740 146.830 125.280 147.000 ;
        RECT 123.740 146.390 125.280 146.560 ;
        RECT 125.450 146.530 125.620 146.860 ;
        RECT 125.950 145.990 127.610 147.400 ;
        RECT 122.890 145.820 127.610 145.990 ;
        RECT 122.890 144.410 123.060 145.820 ;
        RECT 123.400 144.950 123.570 145.280 ;
        RECT 123.740 145.250 125.280 145.420 ;
        RECT 123.740 144.810 125.280 144.980 ;
        RECT 125.450 144.950 125.620 145.280 ;
        RECT 125.950 144.410 127.610 145.820 ;
        RECT 122.890 144.240 127.610 144.410 ;
        RECT 111.540 143.440 111.710 143.790 ;
        RECT 116.680 143.440 116.850 143.790 ;
        RECT 117.190 143.720 122.330 143.890 ;
        RECT 111.925 143.210 116.465 143.380 ;
        RECT 111.540 142.800 111.710 143.150 ;
        RECT 116.680 142.800 116.850 143.150 ;
        RECT 111.925 142.570 116.465 142.740 ;
        RECT 111.540 142.160 111.710 142.510 ;
        RECT 116.680 142.160 116.850 142.510 ;
        RECT 111.925 141.930 116.465 142.100 ;
        RECT 111.540 141.520 111.710 141.870 ;
        RECT 116.680 141.520 116.850 141.870 ;
        RECT 111.925 141.290 116.465 141.460 ;
        RECT 111.540 140.880 111.710 141.230 ;
        RECT 116.680 140.880 116.850 141.230 ;
        RECT 111.925 140.650 116.465 140.820 ;
        RECT 111.540 140.240 111.710 140.590 ;
        RECT 116.680 140.240 116.850 140.590 ;
        RECT 111.925 140.010 116.465 140.180 ;
        RECT 111.540 139.600 111.710 139.950 ;
        RECT 116.680 139.600 116.850 139.950 ;
        RECT 111.925 139.370 116.465 139.540 ;
        RECT 111.540 138.960 111.710 139.310 ;
        RECT 116.680 138.960 116.850 139.310 ;
        RECT 111.925 138.730 116.465 138.900 ;
        RECT 111.540 138.320 111.710 138.670 ;
        RECT 116.680 138.320 116.850 138.670 ;
        RECT 111.925 138.090 116.465 138.260 ;
        RECT 111.540 137.680 111.710 138.030 ;
        RECT 116.680 137.680 116.850 138.030 ;
        RECT 111.925 137.450 116.465 137.620 ;
        RECT 111.540 137.040 111.710 137.390 ;
        RECT 116.680 137.040 116.850 137.390 ;
        RECT 111.925 136.810 116.465 136.980 ;
        RECT 111.540 136.400 111.710 136.750 ;
        RECT 116.680 136.400 116.850 136.750 ;
        RECT 111.925 136.170 116.465 136.340 ;
        RECT 111.540 135.760 111.710 136.110 ;
        RECT 116.680 135.760 116.850 136.110 ;
        RECT 111.925 135.530 116.465 135.700 ;
        RECT 111.540 135.120 111.710 135.470 ;
        RECT 116.680 135.120 116.850 135.470 ;
        RECT 111.925 134.890 116.465 135.060 ;
        RECT 111.540 134.480 111.710 134.830 ;
        RECT 116.680 134.480 116.850 134.830 ;
        RECT 111.925 134.250 116.465 134.420 ;
        RECT 111.540 133.840 111.710 134.190 ;
        RECT 116.680 133.840 116.850 134.190 ;
        RECT 111.925 133.610 116.465 133.780 ;
        RECT 111.540 133.200 111.710 133.550 ;
        RECT 116.680 133.200 116.850 133.550 ;
        RECT 111.925 132.970 116.465 133.140 ;
        RECT 117.190 132.570 118.810 143.720 ;
        RECT 125.950 142.130 127.610 144.240 ;
        RECT 119.490 141.960 127.610 142.130 ;
        RECT 119.490 136.510 119.660 141.960 ;
        RECT 120.340 141.390 124.880 141.560 ;
        RECT 120.000 140.980 120.170 141.330 ;
        RECT 125.050 140.980 125.220 141.330 ;
        RECT 120.340 140.750 124.880 140.920 ;
        RECT 120.000 140.340 120.170 140.690 ;
        RECT 125.050 140.340 125.220 140.690 ;
        RECT 120.340 140.110 124.880 140.280 ;
        RECT 120.000 139.700 120.170 140.050 ;
        RECT 125.050 139.700 125.220 140.050 ;
        RECT 120.340 139.470 124.880 139.640 ;
        RECT 120.000 139.060 120.170 139.410 ;
        RECT 125.050 139.060 125.220 139.410 ;
        RECT 120.340 138.830 124.880 139.000 ;
        RECT 120.000 138.420 120.170 138.770 ;
        RECT 125.050 138.420 125.220 138.770 ;
        RECT 120.340 138.190 124.880 138.360 ;
        RECT 120.000 137.780 120.170 138.130 ;
        RECT 125.050 137.780 125.220 138.130 ;
        RECT 120.340 137.550 124.880 137.720 ;
        RECT 120.000 137.140 120.170 137.490 ;
        RECT 125.050 137.140 125.220 137.490 ;
        RECT 120.340 136.910 124.880 137.080 ;
        RECT 125.560 136.510 127.610 141.960 ;
        RECT 119.490 136.340 127.610 136.510 ;
        RECT 111.030 132.400 118.810 132.570 ;
        RECT 117.190 130.640 118.810 132.400 ;
        RECT 126.410 130.640 127.610 136.340 ;
        RECT 130.290 132.560 130.460 147.840 ;
        RECT 130.940 145.200 131.290 147.360 ;
        RECT 130.940 133.040 131.290 135.200 ;
        RECT 131.770 132.560 131.940 147.840 ;
        RECT 140.200 147.230 142.180 147.920 ;
        RECT 130.290 132.390 131.940 132.560 ;
        RECT 134.040 147.060 142.180 147.230 ;
        RECT 134.040 132.650 134.210 147.060 ;
        RECT 134.935 146.490 139.475 146.660 ;
        RECT 134.550 146.080 134.720 146.430 ;
        RECT 139.690 146.080 139.860 146.430 ;
        RECT 140.200 146.070 142.180 147.060 ;
        RECT 142.515 146.625 142.695 147.445 ;
        RECT 142.905 147.430 144.445 147.600 ;
        RECT 142.905 146.950 144.445 147.120 ;
        RECT 142.905 146.470 144.445 146.640 ;
        RECT 144.655 146.625 144.835 147.445 ;
        RECT 145.170 146.070 145.340 148.000 ;
        RECT 148.960 147.650 150.620 147.920 ;
        RECT 134.935 145.850 139.475 146.020 ;
        RECT 140.200 145.900 145.340 146.070 ;
        RECT 134.550 145.440 134.720 145.790 ;
        RECT 139.690 145.440 139.860 145.790 ;
        RECT 134.935 145.210 139.475 145.380 ;
        RECT 134.550 144.800 134.720 145.150 ;
        RECT 139.690 144.800 139.860 145.150 ;
        RECT 134.935 144.570 139.475 144.740 ;
        RECT 134.550 144.160 134.720 144.510 ;
        RECT 139.690 144.160 139.860 144.510 ;
        RECT 134.935 143.930 139.475 144.100 ;
        RECT 140.200 143.970 142.180 145.900 ;
        RECT 142.515 144.525 142.695 145.345 ;
        RECT 142.905 145.330 144.445 145.500 ;
        RECT 142.905 144.850 144.445 145.020 ;
        RECT 142.905 144.370 144.445 144.540 ;
        RECT 144.655 144.525 144.835 145.345 ;
        RECT 145.170 143.970 145.340 145.900 ;
        RECT 145.900 147.480 150.620 147.650 ;
        RECT 145.900 146.070 146.070 147.480 ;
        RECT 146.410 146.610 146.580 146.940 ;
        RECT 146.750 146.910 148.290 147.080 ;
        RECT 146.750 146.470 148.290 146.640 ;
        RECT 148.460 146.610 148.630 146.940 ;
        RECT 148.960 146.070 150.620 147.480 ;
        RECT 145.900 145.900 150.620 146.070 ;
        RECT 145.900 144.490 146.070 145.900 ;
        RECT 146.410 145.030 146.580 145.360 ;
        RECT 146.750 145.330 148.290 145.500 ;
        RECT 146.750 144.890 148.290 145.060 ;
        RECT 148.460 145.030 148.630 145.360 ;
        RECT 148.960 144.490 150.620 145.900 ;
        RECT 145.900 144.320 150.620 144.490 ;
        RECT 134.550 143.520 134.720 143.870 ;
        RECT 139.690 143.520 139.860 143.870 ;
        RECT 140.200 143.800 145.340 143.970 ;
        RECT 134.935 143.290 139.475 143.460 ;
        RECT 134.550 142.880 134.720 143.230 ;
        RECT 139.690 142.880 139.860 143.230 ;
        RECT 134.935 142.650 139.475 142.820 ;
        RECT 134.550 142.240 134.720 142.590 ;
        RECT 139.690 142.240 139.860 142.590 ;
        RECT 134.935 142.010 139.475 142.180 ;
        RECT 134.550 141.600 134.720 141.950 ;
        RECT 139.690 141.600 139.860 141.950 ;
        RECT 134.935 141.370 139.475 141.540 ;
        RECT 134.550 140.960 134.720 141.310 ;
        RECT 139.690 140.960 139.860 141.310 ;
        RECT 134.935 140.730 139.475 140.900 ;
        RECT 134.550 140.320 134.720 140.670 ;
        RECT 139.690 140.320 139.860 140.670 ;
        RECT 134.935 140.090 139.475 140.260 ;
        RECT 134.550 139.680 134.720 140.030 ;
        RECT 139.690 139.680 139.860 140.030 ;
        RECT 134.935 139.450 139.475 139.620 ;
        RECT 134.550 139.040 134.720 139.390 ;
        RECT 139.690 139.040 139.860 139.390 ;
        RECT 134.935 138.810 139.475 138.980 ;
        RECT 134.550 138.400 134.720 138.750 ;
        RECT 139.690 138.400 139.860 138.750 ;
        RECT 134.935 138.170 139.475 138.340 ;
        RECT 134.550 137.760 134.720 138.110 ;
        RECT 139.690 137.760 139.860 138.110 ;
        RECT 134.935 137.530 139.475 137.700 ;
        RECT 134.550 137.120 134.720 137.470 ;
        RECT 139.690 137.120 139.860 137.470 ;
        RECT 134.935 136.890 139.475 137.060 ;
        RECT 134.550 136.480 134.720 136.830 ;
        RECT 139.690 136.480 139.860 136.830 ;
        RECT 134.935 136.250 139.475 136.420 ;
        RECT 134.550 135.840 134.720 136.190 ;
        RECT 139.690 135.840 139.860 136.190 ;
        RECT 134.935 135.610 139.475 135.780 ;
        RECT 134.550 135.200 134.720 135.550 ;
        RECT 139.690 135.200 139.860 135.550 ;
        RECT 134.935 134.970 139.475 135.140 ;
        RECT 134.550 134.560 134.720 134.910 ;
        RECT 139.690 134.560 139.860 134.910 ;
        RECT 134.935 134.330 139.475 134.500 ;
        RECT 134.550 133.920 134.720 134.270 ;
        RECT 139.690 133.920 139.860 134.270 ;
        RECT 134.935 133.690 139.475 133.860 ;
        RECT 134.550 133.280 134.720 133.630 ;
        RECT 139.690 133.280 139.860 133.630 ;
        RECT 134.935 133.050 139.475 133.220 ;
        RECT 140.200 132.650 141.820 143.800 ;
        RECT 148.960 142.210 150.620 144.320 ;
        RECT 142.500 142.040 150.620 142.210 ;
        RECT 142.500 136.590 142.670 142.040 ;
        RECT 143.350 141.470 147.890 141.640 ;
        RECT 143.010 141.060 143.180 141.410 ;
        RECT 148.060 141.060 148.230 141.410 ;
        RECT 143.350 140.830 147.890 141.000 ;
        RECT 143.010 140.420 143.180 140.770 ;
        RECT 148.060 140.420 148.230 140.770 ;
        RECT 143.350 140.190 147.890 140.360 ;
        RECT 143.010 139.780 143.180 140.130 ;
        RECT 148.060 139.780 148.230 140.130 ;
        RECT 143.350 139.550 147.890 139.720 ;
        RECT 143.010 139.140 143.180 139.490 ;
        RECT 148.060 139.140 148.230 139.490 ;
        RECT 143.350 138.910 147.890 139.080 ;
        RECT 143.010 138.500 143.180 138.850 ;
        RECT 148.060 138.500 148.230 138.850 ;
        RECT 143.350 138.270 147.890 138.440 ;
        RECT 143.010 137.860 143.180 138.210 ;
        RECT 148.060 137.860 148.230 138.210 ;
        RECT 143.350 137.630 147.890 137.800 ;
        RECT 143.010 137.220 143.180 137.570 ;
        RECT 148.060 137.220 148.230 137.570 ;
        RECT 143.350 136.990 147.890 137.160 ;
        RECT 148.570 136.590 150.620 142.040 ;
        RECT 142.500 136.420 150.620 136.590 ;
        RECT 134.040 132.480 141.820 132.650 ;
        RECT 140.200 130.720 141.820 132.480 ;
        RECT 149.420 130.720 150.620 136.420 ;
        RECT 57.730 34.560 60.330 34.730 ;
        RECT 57.730 33.310 57.900 34.560 ;
        RECT 58.530 34.050 59.530 34.220 ;
        RECT 57.730 24.020 57.910 33.310 ;
        RECT 57.730 23.070 57.900 24.020 ;
        RECT 58.300 23.795 58.470 33.835 ;
        RECT 59.590 23.795 59.760 33.835 ;
        RECT 58.530 23.410 59.530 23.580 ;
        RECT 60.160 23.070 60.330 34.560 ;
        RECT 57.730 22.900 60.330 23.070 ;
        RECT 57.680 17.080 60.280 17.250 ;
        RECT 57.680 5.680 57.850 17.080 ;
        RECT 58.480 16.570 59.480 16.740 ;
        RECT 58.250 6.360 58.420 16.400 ;
        RECT 59.540 6.360 59.710 16.400 ;
        RECT 58.480 6.020 59.480 6.190 ;
        RECT 60.110 5.680 60.280 17.080 ;
        RECT 57.680 5.510 60.280 5.680 ;
      LAYER mcon ;
        RECT 61.450 199.440 62.140 199.610 ;
        RECT 61.700 196.875 61.890 198.860 ;
        RECT 61.700 184.720 61.890 186.705 ;
        RECT 65.695 198.080 70.075 198.250 ;
        RECT 65.230 197.750 65.400 197.940 ;
        RECT 70.370 197.750 70.540 197.940 ;
        RECT 65.695 197.440 70.075 197.610 ;
        RECT 65.230 197.110 65.400 197.300 ;
        RECT 70.370 197.110 70.540 197.300 ;
        RECT 65.695 196.800 70.075 196.970 ;
        RECT 65.230 196.470 65.400 196.660 ;
        RECT 70.370 196.470 70.540 196.660 ;
        RECT 65.695 196.160 70.075 196.330 ;
        RECT 65.230 195.830 65.400 196.020 ;
        RECT 70.370 195.830 70.540 196.020 ;
        RECT 65.695 195.520 70.075 195.690 ;
        RECT 65.230 195.190 65.400 195.380 ;
        RECT 70.370 195.190 70.540 195.380 ;
        RECT 65.695 194.880 70.075 195.050 ;
        RECT 65.230 194.550 65.400 194.740 ;
        RECT 70.370 194.550 70.540 194.740 ;
        RECT 65.695 194.240 70.075 194.410 ;
        RECT 65.230 193.910 65.400 194.100 ;
        RECT 70.370 193.910 70.540 194.100 ;
        RECT 65.695 193.600 70.075 193.770 ;
        RECT 65.230 193.270 65.400 193.460 ;
        RECT 70.370 193.270 70.540 193.460 ;
        RECT 65.695 192.960 70.075 193.130 ;
        RECT 65.230 192.630 65.400 192.820 ;
        RECT 70.370 192.630 70.540 192.820 ;
        RECT 65.695 192.320 70.075 192.490 ;
        RECT 65.230 191.990 65.400 192.180 ;
        RECT 70.370 191.990 70.540 192.180 ;
        RECT 65.695 191.680 70.075 191.850 ;
        RECT 65.230 191.350 65.400 191.540 ;
        RECT 70.370 191.350 70.540 191.540 ;
        RECT 65.695 191.040 70.075 191.210 ;
        RECT 65.230 190.710 65.400 190.900 ;
        RECT 70.370 190.710 70.540 190.900 ;
        RECT 65.695 190.400 70.075 190.570 ;
        RECT 65.230 190.070 65.400 190.260 ;
        RECT 70.370 190.070 70.540 190.260 ;
        RECT 65.695 189.760 70.075 189.930 ;
        RECT 65.230 189.430 65.400 189.620 ;
        RECT 70.370 189.430 70.540 189.620 ;
        RECT 65.695 189.120 70.075 189.290 ;
        RECT 65.230 188.790 65.400 188.980 ;
        RECT 70.370 188.790 70.540 188.980 ;
        RECT 65.695 188.480 70.075 188.650 ;
        RECT 65.230 188.150 65.400 188.340 ;
        RECT 70.370 188.150 70.540 188.340 ;
        RECT 65.695 187.840 70.075 188.010 ;
        RECT 65.230 187.510 65.400 187.700 ;
        RECT 70.370 187.510 70.540 187.700 ;
        RECT 65.695 187.200 70.075 187.370 ;
        RECT 65.230 186.870 65.400 187.060 ;
        RECT 70.370 186.870 70.540 187.060 ;
        RECT 65.695 186.560 70.075 186.730 ;
        RECT 65.230 186.230 65.400 186.420 ;
        RECT 70.370 186.230 70.540 186.420 ;
        RECT 65.695 185.920 70.075 186.090 ;
        RECT 65.230 185.590 65.400 185.780 ;
        RECT 70.370 185.590 70.540 185.780 ;
        RECT 65.695 185.280 70.075 185.450 ;
        RECT 65.230 184.950 65.400 185.140 ;
        RECT 70.370 184.950 70.540 185.140 ;
        RECT 65.695 184.640 70.075 184.810 ;
        RECT 71.350 183.710 71.520 199.410 ;
        RECT 72.280 183.710 72.450 199.410 ;
        RECT 73.665 199.020 75.045 199.190 ;
        RECT 73.200 198.780 73.370 198.950 ;
        RECT 75.340 198.780 75.510 198.950 ;
        RECT 73.665 198.540 75.045 198.710 ;
        RECT 73.200 198.300 73.370 198.470 ;
        RECT 75.340 198.300 75.510 198.470 ;
        RECT 73.665 198.060 75.045 198.230 ;
        RECT 73.665 196.920 75.045 197.090 ;
        RECT 73.200 196.680 73.370 196.850 ;
        RECT 75.340 196.680 75.510 196.850 ;
        RECT 73.665 196.440 75.045 196.610 ;
        RECT 73.200 196.200 73.370 196.370 ;
        RECT 75.340 196.200 75.510 196.370 ;
        RECT 73.665 195.960 75.045 196.130 ;
        RECT 77.510 198.500 78.890 198.670 ;
        RECT 77.090 198.280 77.260 198.450 ;
        RECT 79.140 198.280 79.310 198.450 ;
        RECT 77.510 198.060 78.890 198.230 ;
        RECT 80.200 198.410 81.200 199.410 ;
        RECT 77.510 196.920 78.890 197.090 ;
        RECT 77.090 196.700 77.260 196.870 ;
        RECT 79.140 196.700 79.310 196.870 ;
        RECT 77.510 196.480 78.890 196.650 ;
        RECT 74.110 193.060 78.490 193.230 ;
        RECT 73.690 192.730 73.860 192.920 ;
        RECT 78.740 192.730 78.910 192.920 ;
        RECT 74.110 192.420 78.490 192.590 ;
        RECT 73.690 192.090 73.860 192.280 ;
        RECT 78.740 192.090 78.910 192.280 ;
        RECT 74.110 191.780 78.490 191.950 ;
        RECT 73.690 191.450 73.860 191.640 ;
        RECT 78.740 191.450 78.910 191.640 ;
        RECT 74.110 191.140 78.490 191.310 ;
        RECT 73.690 190.810 73.860 191.000 ;
        RECT 78.740 190.810 78.910 191.000 ;
        RECT 74.110 190.500 78.490 190.670 ;
        RECT 73.690 190.170 73.860 190.360 ;
        RECT 78.740 190.170 78.910 190.360 ;
        RECT 74.110 189.860 78.490 190.030 ;
        RECT 73.690 189.530 73.860 189.720 ;
        RECT 78.740 189.530 78.910 189.720 ;
        RECT 74.110 189.220 78.490 189.390 ;
        RECT 73.690 188.890 73.860 189.080 ;
        RECT 78.740 188.890 78.910 189.080 ;
        RECT 74.110 188.580 78.490 188.750 ;
        RECT 71.400 182.410 72.400 183.410 ;
        RECT 80.150 182.410 80.320 198.110 ;
        RECT 86.190 199.360 86.880 199.530 ;
        RECT 86.440 196.795 86.630 198.780 ;
        RECT 86.440 184.640 86.630 186.625 ;
        RECT 90.435 198.000 94.815 198.170 ;
        RECT 89.970 197.670 90.140 197.860 ;
        RECT 95.110 197.670 95.280 197.860 ;
        RECT 90.435 197.360 94.815 197.530 ;
        RECT 89.970 197.030 90.140 197.220 ;
        RECT 95.110 197.030 95.280 197.220 ;
        RECT 90.435 196.720 94.815 196.890 ;
        RECT 89.970 196.390 90.140 196.580 ;
        RECT 95.110 196.390 95.280 196.580 ;
        RECT 90.435 196.080 94.815 196.250 ;
        RECT 89.970 195.750 90.140 195.940 ;
        RECT 95.110 195.750 95.280 195.940 ;
        RECT 90.435 195.440 94.815 195.610 ;
        RECT 89.970 195.110 90.140 195.300 ;
        RECT 95.110 195.110 95.280 195.300 ;
        RECT 90.435 194.800 94.815 194.970 ;
        RECT 89.970 194.470 90.140 194.660 ;
        RECT 95.110 194.470 95.280 194.660 ;
        RECT 90.435 194.160 94.815 194.330 ;
        RECT 89.970 193.830 90.140 194.020 ;
        RECT 95.110 193.830 95.280 194.020 ;
        RECT 90.435 193.520 94.815 193.690 ;
        RECT 89.970 193.190 90.140 193.380 ;
        RECT 95.110 193.190 95.280 193.380 ;
        RECT 90.435 192.880 94.815 193.050 ;
        RECT 89.970 192.550 90.140 192.740 ;
        RECT 95.110 192.550 95.280 192.740 ;
        RECT 90.435 192.240 94.815 192.410 ;
        RECT 89.970 191.910 90.140 192.100 ;
        RECT 95.110 191.910 95.280 192.100 ;
        RECT 90.435 191.600 94.815 191.770 ;
        RECT 89.970 191.270 90.140 191.460 ;
        RECT 95.110 191.270 95.280 191.460 ;
        RECT 90.435 190.960 94.815 191.130 ;
        RECT 89.970 190.630 90.140 190.820 ;
        RECT 95.110 190.630 95.280 190.820 ;
        RECT 90.435 190.320 94.815 190.490 ;
        RECT 89.970 189.990 90.140 190.180 ;
        RECT 95.110 189.990 95.280 190.180 ;
        RECT 90.435 189.680 94.815 189.850 ;
        RECT 89.970 189.350 90.140 189.540 ;
        RECT 95.110 189.350 95.280 189.540 ;
        RECT 90.435 189.040 94.815 189.210 ;
        RECT 89.970 188.710 90.140 188.900 ;
        RECT 95.110 188.710 95.280 188.900 ;
        RECT 90.435 188.400 94.815 188.570 ;
        RECT 89.970 188.070 90.140 188.260 ;
        RECT 95.110 188.070 95.280 188.260 ;
        RECT 90.435 187.760 94.815 187.930 ;
        RECT 89.970 187.430 90.140 187.620 ;
        RECT 95.110 187.430 95.280 187.620 ;
        RECT 90.435 187.120 94.815 187.290 ;
        RECT 89.970 186.790 90.140 186.980 ;
        RECT 95.110 186.790 95.280 186.980 ;
        RECT 90.435 186.480 94.815 186.650 ;
        RECT 89.970 186.150 90.140 186.340 ;
        RECT 95.110 186.150 95.280 186.340 ;
        RECT 90.435 185.840 94.815 186.010 ;
        RECT 89.970 185.510 90.140 185.700 ;
        RECT 95.110 185.510 95.280 185.700 ;
        RECT 90.435 185.200 94.815 185.370 ;
        RECT 89.970 184.870 90.140 185.060 ;
        RECT 95.110 184.870 95.280 185.060 ;
        RECT 90.435 184.560 94.815 184.730 ;
        RECT 96.090 183.630 96.260 199.330 ;
        RECT 97.020 183.630 97.190 199.330 ;
        RECT 98.405 198.940 99.785 199.110 ;
        RECT 97.940 198.700 98.110 198.870 ;
        RECT 100.080 198.700 100.250 198.870 ;
        RECT 98.405 198.460 99.785 198.630 ;
        RECT 97.940 198.220 98.110 198.390 ;
        RECT 100.080 198.220 100.250 198.390 ;
        RECT 98.405 197.980 99.785 198.150 ;
        RECT 98.405 196.840 99.785 197.010 ;
        RECT 97.940 196.600 98.110 196.770 ;
        RECT 100.080 196.600 100.250 196.770 ;
        RECT 98.405 196.360 99.785 196.530 ;
        RECT 97.940 196.120 98.110 196.290 ;
        RECT 100.080 196.120 100.250 196.290 ;
        RECT 98.405 195.880 99.785 196.050 ;
        RECT 102.250 198.420 103.630 198.590 ;
        RECT 101.830 198.200 102.000 198.370 ;
        RECT 103.880 198.200 104.050 198.370 ;
        RECT 102.250 197.980 103.630 198.150 ;
        RECT 104.940 198.330 105.940 199.330 ;
        RECT 102.250 196.840 103.630 197.010 ;
        RECT 101.830 196.620 102.000 196.790 ;
        RECT 103.880 196.620 104.050 196.790 ;
        RECT 102.250 196.400 103.630 196.570 ;
        RECT 98.850 192.980 103.230 193.150 ;
        RECT 98.430 192.650 98.600 192.840 ;
        RECT 103.480 192.650 103.650 192.840 ;
        RECT 98.850 192.340 103.230 192.510 ;
        RECT 98.430 192.010 98.600 192.200 ;
        RECT 103.480 192.010 103.650 192.200 ;
        RECT 98.850 191.700 103.230 191.870 ;
        RECT 98.430 191.370 98.600 191.560 ;
        RECT 103.480 191.370 103.650 191.560 ;
        RECT 98.850 191.060 103.230 191.230 ;
        RECT 98.430 190.730 98.600 190.920 ;
        RECT 103.480 190.730 103.650 190.920 ;
        RECT 98.850 190.420 103.230 190.590 ;
        RECT 98.430 190.090 98.600 190.280 ;
        RECT 103.480 190.090 103.650 190.280 ;
        RECT 98.850 189.780 103.230 189.950 ;
        RECT 98.430 189.450 98.600 189.640 ;
        RECT 103.480 189.450 103.650 189.640 ;
        RECT 98.850 189.140 103.230 189.310 ;
        RECT 98.430 188.810 98.600 189.000 ;
        RECT 103.480 188.810 103.650 189.000 ;
        RECT 98.850 188.500 103.230 188.670 ;
        RECT 96.140 182.330 97.140 183.330 ;
        RECT 104.890 182.330 105.060 198.030 ;
        RECT 109.440 199.350 110.130 199.520 ;
        RECT 109.690 196.785 109.880 198.770 ;
        RECT 109.690 184.630 109.880 186.615 ;
        RECT 113.685 197.990 118.065 198.160 ;
        RECT 113.220 197.660 113.390 197.850 ;
        RECT 118.360 197.660 118.530 197.850 ;
        RECT 113.685 197.350 118.065 197.520 ;
        RECT 113.220 197.020 113.390 197.210 ;
        RECT 118.360 197.020 118.530 197.210 ;
        RECT 113.685 196.710 118.065 196.880 ;
        RECT 113.220 196.380 113.390 196.570 ;
        RECT 118.360 196.380 118.530 196.570 ;
        RECT 113.685 196.070 118.065 196.240 ;
        RECT 113.220 195.740 113.390 195.930 ;
        RECT 118.360 195.740 118.530 195.930 ;
        RECT 113.685 195.430 118.065 195.600 ;
        RECT 113.220 195.100 113.390 195.290 ;
        RECT 118.360 195.100 118.530 195.290 ;
        RECT 113.685 194.790 118.065 194.960 ;
        RECT 113.220 194.460 113.390 194.650 ;
        RECT 118.360 194.460 118.530 194.650 ;
        RECT 113.685 194.150 118.065 194.320 ;
        RECT 113.220 193.820 113.390 194.010 ;
        RECT 118.360 193.820 118.530 194.010 ;
        RECT 113.685 193.510 118.065 193.680 ;
        RECT 113.220 193.180 113.390 193.370 ;
        RECT 118.360 193.180 118.530 193.370 ;
        RECT 113.685 192.870 118.065 193.040 ;
        RECT 113.220 192.540 113.390 192.730 ;
        RECT 118.360 192.540 118.530 192.730 ;
        RECT 113.685 192.230 118.065 192.400 ;
        RECT 113.220 191.900 113.390 192.090 ;
        RECT 118.360 191.900 118.530 192.090 ;
        RECT 113.685 191.590 118.065 191.760 ;
        RECT 113.220 191.260 113.390 191.450 ;
        RECT 118.360 191.260 118.530 191.450 ;
        RECT 113.685 190.950 118.065 191.120 ;
        RECT 113.220 190.620 113.390 190.810 ;
        RECT 118.360 190.620 118.530 190.810 ;
        RECT 113.685 190.310 118.065 190.480 ;
        RECT 113.220 189.980 113.390 190.170 ;
        RECT 118.360 189.980 118.530 190.170 ;
        RECT 113.685 189.670 118.065 189.840 ;
        RECT 113.220 189.340 113.390 189.530 ;
        RECT 118.360 189.340 118.530 189.530 ;
        RECT 113.685 189.030 118.065 189.200 ;
        RECT 113.220 188.700 113.390 188.890 ;
        RECT 118.360 188.700 118.530 188.890 ;
        RECT 113.685 188.390 118.065 188.560 ;
        RECT 113.220 188.060 113.390 188.250 ;
        RECT 118.360 188.060 118.530 188.250 ;
        RECT 113.685 187.750 118.065 187.920 ;
        RECT 113.220 187.420 113.390 187.610 ;
        RECT 118.360 187.420 118.530 187.610 ;
        RECT 113.685 187.110 118.065 187.280 ;
        RECT 113.220 186.780 113.390 186.970 ;
        RECT 118.360 186.780 118.530 186.970 ;
        RECT 113.685 186.470 118.065 186.640 ;
        RECT 113.220 186.140 113.390 186.330 ;
        RECT 118.360 186.140 118.530 186.330 ;
        RECT 113.685 185.830 118.065 186.000 ;
        RECT 113.220 185.500 113.390 185.690 ;
        RECT 118.360 185.500 118.530 185.690 ;
        RECT 113.685 185.190 118.065 185.360 ;
        RECT 113.220 184.860 113.390 185.050 ;
        RECT 118.360 184.860 118.530 185.050 ;
        RECT 113.685 184.550 118.065 184.720 ;
        RECT 119.340 183.620 119.510 199.320 ;
        RECT 120.270 183.620 120.440 199.320 ;
        RECT 121.655 198.930 123.035 199.100 ;
        RECT 121.190 198.690 121.360 198.860 ;
        RECT 123.330 198.690 123.500 198.860 ;
        RECT 121.655 198.450 123.035 198.620 ;
        RECT 121.190 198.210 121.360 198.380 ;
        RECT 123.330 198.210 123.500 198.380 ;
        RECT 121.655 197.970 123.035 198.140 ;
        RECT 121.655 196.830 123.035 197.000 ;
        RECT 121.190 196.590 121.360 196.760 ;
        RECT 123.330 196.590 123.500 196.760 ;
        RECT 121.655 196.350 123.035 196.520 ;
        RECT 121.190 196.110 121.360 196.280 ;
        RECT 123.330 196.110 123.500 196.280 ;
        RECT 121.655 195.870 123.035 196.040 ;
        RECT 125.500 198.410 126.880 198.580 ;
        RECT 125.080 198.190 125.250 198.360 ;
        RECT 127.130 198.190 127.300 198.360 ;
        RECT 125.500 197.970 126.880 198.140 ;
        RECT 128.190 198.320 129.190 199.320 ;
        RECT 125.500 196.830 126.880 197.000 ;
        RECT 125.080 196.610 125.250 196.780 ;
        RECT 127.130 196.610 127.300 196.780 ;
        RECT 125.500 196.390 126.880 196.560 ;
        RECT 122.100 192.970 126.480 193.140 ;
        RECT 121.680 192.640 121.850 192.830 ;
        RECT 126.730 192.640 126.900 192.830 ;
        RECT 122.100 192.330 126.480 192.500 ;
        RECT 121.680 192.000 121.850 192.190 ;
        RECT 126.730 192.000 126.900 192.190 ;
        RECT 122.100 191.690 126.480 191.860 ;
        RECT 121.680 191.360 121.850 191.550 ;
        RECT 126.730 191.360 126.900 191.550 ;
        RECT 122.100 191.050 126.480 191.220 ;
        RECT 121.680 190.720 121.850 190.910 ;
        RECT 126.730 190.720 126.900 190.910 ;
        RECT 122.100 190.410 126.480 190.580 ;
        RECT 121.680 190.080 121.850 190.270 ;
        RECT 126.730 190.080 126.900 190.270 ;
        RECT 122.100 189.770 126.480 189.940 ;
        RECT 121.680 189.440 121.850 189.630 ;
        RECT 126.730 189.440 126.900 189.630 ;
        RECT 122.100 189.130 126.480 189.300 ;
        RECT 121.680 188.800 121.850 188.990 ;
        RECT 126.730 188.800 126.900 188.990 ;
        RECT 122.100 188.490 126.480 188.660 ;
        RECT 119.390 182.320 120.390 183.320 ;
        RECT 128.140 182.320 128.310 198.020 ;
        RECT 133.070 199.340 133.760 199.510 ;
        RECT 133.320 196.775 133.510 198.760 ;
        RECT 133.320 184.620 133.510 186.605 ;
        RECT 137.315 197.980 141.695 198.150 ;
        RECT 136.850 197.650 137.020 197.840 ;
        RECT 141.990 197.650 142.160 197.840 ;
        RECT 137.315 197.340 141.695 197.510 ;
        RECT 136.850 197.010 137.020 197.200 ;
        RECT 141.990 197.010 142.160 197.200 ;
        RECT 137.315 196.700 141.695 196.870 ;
        RECT 136.850 196.370 137.020 196.560 ;
        RECT 141.990 196.370 142.160 196.560 ;
        RECT 137.315 196.060 141.695 196.230 ;
        RECT 136.850 195.730 137.020 195.920 ;
        RECT 141.990 195.730 142.160 195.920 ;
        RECT 137.315 195.420 141.695 195.590 ;
        RECT 136.850 195.090 137.020 195.280 ;
        RECT 141.990 195.090 142.160 195.280 ;
        RECT 137.315 194.780 141.695 194.950 ;
        RECT 136.850 194.450 137.020 194.640 ;
        RECT 141.990 194.450 142.160 194.640 ;
        RECT 137.315 194.140 141.695 194.310 ;
        RECT 136.850 193.810 137.020 194.000 ;
        RECT 141.990 193.810 142.160 194.000 ;
        RECT 137.315 193.500 141.695 193.670 ;
        RECT 136.850 193.170 137.020 193.360 ;
        RECT 141.990 193.170 142.160 193.360 ;
        RECT 137.315 192.860 141.695 193.030 ;
        RECT 136.850 192.530 137.020 192.720 ;
        RECT 141.990 192.530 142.160 192.720 ;
        RECT 137.315 192.220 141.695 192.390 ;
        RECT 136.850 191.890 137.020 192.080 ;
        RECT 141.990 191.890 142.160 192.080 ;
        RECT 137.315 191.580 141.695 191.750 ;
        RECT 136.850 191.250 137.020 191.440 ;
        RECT 141.990 191.250 142.160 191.440 ;
        RECT 137.315 190.940 141.695 191.110 ;
        RECT 136.850 190.610 137.020 190.800 ;
        RECT 141.990 190.610 142.160 190.800 ;
        RECT 137.315 190.300 141.695 190.470 ;
        RECT 136.850 189.970 137.020 190.160 ;
        RECT 141.990 189.970 142.160 190.160 ;
        RECT 137.315 189.660 141.695 189.830 ;
        RECT 136.850 189.330 137.020 189.520 ;
        RECT 141.990 189.330 142.160 189.520 ;
        RECT 137.315 189.020 141.695 189.190 ;
        RECT 136.850 188.690 137.020 188.880 ;
        RECT 141.990 188.690 142.160 188.880 ;
        RECT 137.315 188.380 141.695 188.550 ;
        RECT 136.850 188.050 137.020 188.240 ;
        RECT 141.990 188.050 142.160 188.240 ;
        RECT 137.315 187.740 141.695 187.910 ;
        RECT 136.850 187.410 137.020 187.600 ;
        RECT 141.990 187.410 142.160 187.600 ;
        RECT 137.315 187.100 141.695 187.270 ;
        RECT 136.850 186.770 137.020 186.960 ;
        RECT 141.990 186.770 142.160 186.960 ;
        RECT 137.315 186.460 141.695 186.630 ;
        RECT 136.850 186.130 137.020 186.320 ;
        RECT 141.990 186.130 142.160 186.320 ;
        RECT 137.315 185.820 141.695 185.990 ;
        RECT 136.850 185.490 137.020 185.680 ;
        RECT 141.990 185.490 142.160 185.680 ;
        RECT 137.315 185.180 141.695 185.350 ;
        RECT 136.850 184.850 137.020 185.040 ;
        RECT 141.990 184.850 142.160 185.040 ;
        RECT 137.315 184.540 141.695 184.710 ;
        RECT 142.970 183.610 143.140 199.310 ;
        RECT 143.900 183.610 144.070 199.310 ;
        RECT 145.285 198.920 146.665 199.090 ;
        RECT 144.820 198.680 144.990 198.850 ;
        RECT 146.960 198.680 147.130 198.850 ;
        RECT 145.285 198.440 146.665 198.610 ;
        RECT 144.820 198.200 144.990 198.370 ;
        RECT 146.960 198.200 147.130 198.370 ;
        RECT 145.285 197.960 146.665 198.130 ;
        RECT 145.285 196.820 146.665 196.990 ;
        RECT 144.820 196.580 144.990 196.750 ;
        RECT 146.960 196.580 147.130 196.750 ;
        RECT 145.285 196.340 146.665 196.510 ;
        RECT 144.820 196.100 144.990 196.270 ;
        RECT 146.960 196.100 147.130 196.270 ;
        RECT 145.285 195.860 146.665 196.030 ;
        RECT 149.130 198.400 150.510 198.570 ;
        RECT 148.710 198.180 148.880 198.350 ;
        RECT 150.760 198.180 150.930 198.350 ;
        RECT 149.130 197.960 150.510 198.130 ;
        RECT 151.820 198.310 152.820 199.310 ;
        RECT 149.130 196.820 150.510 196.990 ;
        RECT 148.710 196.600 148.880 196.770 ;
        RECT 150.760 196.600 150.930 196.770 ;
        RECT 149.130 196.380 150.510 196.550 ;
        RECT 145.730 192.960 150.110 193.130 ;
        RECT 145.310 192.630 145.480 192.820 ;
        RECT 150.360 192.630 150.530 192.820 ;
        RECT 145.730 192.320 150.110 192.490 ;
        RECT 145.310 191.990 145.480 192.180 ;
        RECT 150.360 191.990 150.530 192.180 ;
        RECT 145.730 191.680 150.110 191.850 ;
        RECT 145.310 191.350 145.480 191.540 ;
        RECT 150.360 191.350 150.530 191.540 ;
        RECT 145.730 191.040 150.110 191.210 ;
        RECT 145.310 190.710 145.480 190.900 ;
        RECT 150.360 190.710 150.530 190.900 ;
        RECT 145.730 190.400 150.110 190.570 ;
        RECT 145.310 190.070 145.480 190.260 ;
        RECT 150.360 190.070 150.530 190.260 ;
        RECT 145.730 189.760 150.110 189.930 ;
        RECT 145.310 189.430 145.480 189.620 ;
        RECT 150.360 189.430 150.530 189.620 ;
        RECT 145.730 189.120 150.110 189.290 ;
        RECT 145.310 188.790 145.480 188.980 ;
        RECT 150.360 188.790 150.530 188.980 ;
        RECT 145.730 188.480 150.110 188.650 ;
        RECT 143.020 182.310 144.020 183.310 ;
        RECT 151.770 182.310 151.940 198.010 ;
        RECT 61.340 173.350 62.030 173.520 ;
        RECT 61.590 170.785 61.780 172.770 ;
        RECT 61.590 158.630 61.780 160.615 ;
        RECT 65.585 171.990 69.965 172.160 ;
        RECT 65.120 171.660 65.290 171.850 ;
        RECT 70.260 171.660 70.430 171.850 ;
        RECT 65.585 171.350 69.965 171.520 ;
        RECT 65.120 171.020 65.290 171.210 ;
        RECT 70.260 171.020 70.430 171.210 ;
        RECT 65.585 170.710 69.965 170.880 ;
        RECT 65.120 170.380 65.290 170.570 ;
        RECT 70.260 170.380 70.430 170.570 ;
        RECT 65.585 170.070 69.965 170.240 ;
        RECT 65.120 169.740 65.290 169.930 ;
        RECT 70.260 169.740 70.430 169.930 ;
        RECT 65.585 169.430 69.965 169.600 ;
        RECT 65.120 169.100 65.290 169.290 ;
        RECT 70.260 169.100 70.430 169.290 ;
        RECT 65.585 168.790 69.965 168.960 ;
        RECT 65.120 168.460 65.290 168.650 ;
        RECT 70.260 168.460 70.430 168.650 ;
        RECT 65.585 168.150 69.965 168.320 ;
        RECT 65.120 167.820 65.290 168.010 ;
        RECT 70.260 167.820 70.430 168.010 ;
        RECT 65.585 167.510 69.965 167.680 ;
        RECT 65.120 167.180 65.290 167.370 ;
        RECT 70.260 167.180 70.430 167.370 ;
        RECT 65.585 166.870 69.965 167.040 ;
        RECT 65.120 166.540 65.290 166.730 ;
        RECT 70.260 166.540 70.430 166.730 ;
        RECT 65.585 166.230 69.965 166.400 ;
        RECT 65.120 165.900 65.290 166.090 ;
        RECT 70.260 165.900 70.430 166.090 ;
        RECT 65.585 165.590 69.965 165.760 ;
        RECT 65.120 165.260 65.290 165.450 ;
        RECT 70.260 165.260 70.430 165.450 ;
        RECT 65.585 164.950 69.965 165.120 ;
        RECT 65.120 164.620 65.290 164.810 ;
        RECT 70.260 164.620 70.430 164.810 ;
        RECT 65.585 164.310 69.965 164.480 ;
        RECT 65.120 163.980 65.290 164.170 ;
        RECT 70.260 163.980 70.430 164.170 ;
        RECT 65.585 163.670 69.965 163.840 ;
        RECT 65.120 163.340 65.290 163.530 ;
        RECT 70.260 163.340 70.430 163.530 ;
        RECT 65.585 163.030 69.965 163.200 ;
        RECT 65.120 162.700 65.290 162.890 ;
        RECT 70.260 162.700 70.430 162.890 ;
        RECT 65.585 162.390 69.965 162.560 ;
        RECT 65.120 162.060 65.290 162.250 ;
        RECT 70.260 162.060 70.430 162.250 ;
        RECT 65.585 161.750 69.965 161.920 ;
        RECT 65.120 161.420 65.290 161.610 ;
        RECT 70.260 161.420 70.430 161.610 ;
        RECT 65.585 161.110 69.965 161.280 ;
        RECT 65.120 160.780 65.290 160.970 ;
        RECT 70.260 160.780 70.430 160.970 ;
        RECT 65.585 160.470 69.965 160.640 ;
        RECT 65.120 160.140 65.290 160.330 ;
        RECT 70.260 160.140 70.430 160.330 ;
        RECT 65.585 159.830 69.965 160.000 ;
        RECT 65.120 159.500 65.290 159.690 ;
        RECT 70.260 159.500 70.430 159.690 ;
        RECT 65.585 159.190 69.965 159.360 ;
        RECT 65.120 158.860 65.290 159.050 ;
        RECT 70.260 158.860 70.430 159.050 ;
        RECT 65.585 158.550 69.965 158.720 ;
        RECT 71.240 157.620 71.410 173.320 ;
        RECT 72.170 157.620 72.340 173.320 ;
        RECT 73.555 172.930 74.935 173.100 ;
        RECT 73.090 172.690 73.260 172.860 ;
        RECT 75.230 172.690 75.400 172.860 ;
        RECT 73.555 172.450 74.935 172.620 ;
        RECT 73.090 172.210 73.260 172.380 ;
        RECT 75.230 172.210 75.400 172.380 ;
        RECT 73.555 171.970 74.935 172.140 ;
        RECT 73.555 170.830 74.935 171.000 ;
        RECT 73.090 170.590 73.260 170.760 ;
        RECT 75.230 170.590 75.400 170.760 ;
        RECT 73.555 170.350 74.935 170.520 ;
        RECT 73.090 170.110 73.260 170.280 ;
        RECT 75.230 170.110 75.400 170.280 ;
        RECT 73.555 169.870 74.935 170.040 ;
        RECT 77.400 172.410 78.780 172.580 ;
        RECT 76.980 172.190 77.150 172.360 ;
        RECT 79.030 172.190 79.200 172.360 ;
        RECT 77.400 171.970 78.780 172.140 ;
        RECT 80.090 172.320 81.090 173.320 ;
        RECT 77.400 170.830 78.780 171.000 ;
        RECT 76.980 170.610 77.150 170.780 ;
        RECT 79.030 170.610 79.200 170.780 ;
        RECT 77.400 170.390 78.780 170.560 ;
        RECT 74.000 166.970 78.380 167.140 ;
        RECT 73.580 166.640 73.750 166.830 ;
        RECT 78.630 166.640 78.800 166.830 ;
        RECT 74.000 166.330 78.380 166.500 ;
        RECT 73.580 166.000 73.750 166.190 ;
        RECT 78.630 166.000 78.800 166.190 ;
        RECT 74.000 165.690 78.380 165.860 ;
        RECT 73.580 165.360 73.750 165.550 ;
        RECT 78.630 165.360 78.800 165.550 ;
        RECT 74.000 165.050 78.380 165.220 ;
        RECT 73.580 164.720 73.750 164.910 ;
        RECT 78.630 164.720 78.800 164.910 ;
        RECT 74.000 164.410 78.380 164.580 ;
        RECT 73.580 164.080 73.750 164.270 ;
        RECT 78.630 164.080 78.800 164.270 ;
        RECT 74.000 163.770 78.380 163.940 ;
        RECT 73.580 163.440 73.750 163.630 ;
        RECT 78.630 163.440 78.800 163.630 ;
        RECT 74.000 163.130 78.380 163.300 ;
        RECT 73.580 162.800 73.750 162.990 ;
        RECT 78.630 162.800 78.800 162.990 ;
        RECT 74.000 162.490 78.380 162.660 ;
        RECT 71.290 156.320 72.290 157.320 ;
        RECT 80.040 156.320 80.210 172.020 ;
        RECT 84.520 173.260 85.210 173.430 ;
        RECT 84.770 170.695 84.960 172.680 ;
        RECT 84.770 158.540 84.960 160.525 ;
        RECT 88.765 171.900 93.145 172.070 ;
        RECT 88.300 171.570 88.470 171.760 ;
        RECT 93.440 171.570 93.610 171.760 ;
        RECT 88.765 171.260 93.145 171.430 ;
        RECT 88.300 170.930 88.470 171.120 ;
        RECT 93.440 170.930 93.610 171.120 ;
        RECT 88.765 170.620 93.145 170.790 ;
        RECT 88.300 170.290 88.470 170.480 ;
        RECT 93.440 170.290 93.610 170.480 ;
        RECT 88.765 169.980 93.145 170.150 ;
        RECT 88.300 169.650 88.470 169.840 ;
        RECT 93.440 169.650 93.610 169.840 ;
        RECT 88.765 169.340 93.145 169.510 ;
        RECT 88.300 169.010 88.470 169.200 ;
        RECT 93.440 169.010 93.610 169.200 ;
        RECT 88.765 168.700 93.145 168.870 ;
        RECT 88.300 168.370 88.470 168.560 ;
        RECT 93.440 168.370 93.610 168.560 ;
        RECT 88.765 168.060 93.145 168.230 ;
        RECT 88.300 167.730 88.470 167.920 ;
        RECT 93.440 167.730 93.610 167.920 ;
        RECT 88.765 167.420 93.145 167.590 ;
        RECT 88.300 167.090 88.470 167.280 ;
        RECT 93.440 167.090 93.610 167.280 ;
        RECT 88.765 166.780 93.145 166.950 ;
        RECT 88.300 166.450 88.470 166.640 ;
        RECT 93.440 166.450 93.610 166.640 ;
        RECT 88.765 166.140 93.145 166.310 ;
        RECT 88.300 165.810 88.470 166.000 ;
        RECT 93.440 165.810 93.610 166.000 ;
        RECT 88.765 165.500 93.145 165.670 ;
        RECT 88.300 165.170 88.470 165.360 ;
        RECT 93.440 165.170 93.610 165.360 ;
        RECT 88.765 164.860 93.145 165.030 ;
        RECT 88.300 164.530 88.470 164.720 ;
        RECT 93.440 164.530 93.610 164.720 ;
        RECT 88.765 164.220 93.145 164.390 ;
        RECT 88.300 163.890 88.470 164.080 ;
        RECT 93.440 163.890 93.610 164.080 ;
        RECT 88.765 163.580 93.145 163.750 ;
        RECT 88.300 163.250 88.470 163.440 ;
        RECT 93.440 163.250 93.610 163.440 ;
        RECT 88.765 162.940 93.145 163.110 ;
        RECT 88.300 162.610 88.470 162.800 ;
        RECT 93.440 162.610 93.610 162.800 ;
        RECT 88.765 162.300 93.145 162.470 ;
        RECT 88.300 161.970 88.470 162.160 ;
        RECT 93.440 161.970 93.610 162.160 ;
        RECT 88.765 161.660 93.145 161.830 ;
        RECT 88.300 161.330 88.470 161.520 ;
        RECT 93.440 161.330 93.610 161.520 ;
        RECT 88.765 161.020 93.145 161.190 ;
        RECT 88.300 160.690 88.470 160.880 ;
        RECT 93.440 160.690 93.610 160.880 ;
        RECT 88.765 160.380 93.145 160.550 ;
        RECT 88.300 160.050 88.470 160.240 ;
        RECT 93.440 160.050 93.610 160.240 ;
        RECT 88.765 159.740 93.145 159.910 ;
        RECT 88.300 159.410 88.470 159.600 ;
        RECT 93.440 159.410 93.610 159.600 ;
        RECT 88.765 159.100 93.145 159.270 ;
        RECT 88.300 158.770 88.470 158.960 ;
        RECT 93.440 158.770 93.610 158.960 ;
        RECT 88.765 158.460 93.145 158.630 ;
        RECT 94.420 157.530 94.590 173.230 ;
        RECT 95.350 157.530 95.520 173.230 ;
        RECT 96.735 172.840 98.115 173.010 ;
        RECT 96.270 172.600 96.440 172.770 ;
        RECT 98.410 172.600 98.580 172.770 ;
        RECT 96.735 172.360 98.115 172.530 ;
        RECT 96.270 172.120 96.440 172.290 ;
        RECT 98.410 172.120 98.580 172.290 ;
        RECT 96.735 171.880 98.115 172.050 ;
        RECT 107.420 173.460 108.110 173.630 ;
        RECT 96.735 170.740 98.115 170.910 ;
        RECT 96.270 170.500 96.440 170.670 ;
        RECT 98.410 170.500 98.580 170.670 ;
        RECT 96.735 170.260 98.115 170.430 ;
        RECT 96.270 170.020 96.440 170.190 ;
        RECT 98.410 170.020 98.580 170.190 ;
        RECT 96.735 169.780 98.115 169.950 ;
        RECT 100.580 172.320 101.960 172.490 ;
        RECT 100.160 172.100 100.330 172.270 ;
        RECT 102.210 172.100 102.380 172.270 ;
        RECT 100.580 171.880 101.960 172.050 ;
        RECT 103.270 172.230 104.270 173.230 ;
        RECT 100.580 170.740 101.960 170.910 ;
        RECT 100.160 170.520 100.330 170.690 ;
        RECT 102.210 170.520 102.380 170.690 ;
        RECT 100.580 170.300 101.960 170.470 ;
        RECT 97.180 166.880 101.560 167.050 ;
        RECT 96.760 166.550 96.930 166.740 ;
        RECT 101.810 166.550 101.980 166.740 ;
        RECT 97.180 166.240 101.560 166.410 ;
        RECT 96.760 165.910 96.930 166.100 ;
        RECT 101.810 165.910 101.980 166.100 ;
        RECT 97.180 165.600 101.560 165.770 ;
        RECT 96.760 165.270 96.930 165.460 ;
        RECT 101.810 165.270 101.980 165.460 ;
        RECT 97.180 164.960 101.560 165.130 ;
        RECT 96.760 164.630 96.930 164.820 ;
        RECT 101.810 164.630 101.980 164.820 ;
        RECT 97.180 164.320 101.560 164.490 ;
        RECT 96.760 163.990 96.930 164.180 ;
        RECT 101.810 163.990 101.980 164.180 ;
        RECT 97.180 163.680 101.560 163.850 ;
        RECT 96.760 163.350 96.930 163.540 ;
        RECT 101.810 163.350 101.980 163.540 ;
        RECT 97.180 163.040 101.560 163.210 ;
        RECT 96.760 162.710 96.930 162.900 ;
        RECT 101.810 162.710 101.980 162.900 ;
        RECT 97.180 162.400 101.560 162.570 ;
        RECT 94.470 156.230 95.470 157.230 ;
        RECT 103.220 156.230 103.390 171.930 ;
        RECT 107.670 170.895 107.860 172.880 ;
        RECT 107.670 158.740 107.860 160.725 ;
        RECT 111.665 172.100 116.045 172.270 ;
        RECT 111.200 171.770 111.370 171.960 ;
        RECT 116.340 171.770 116.510 171.960 ;
        RECT 111.665 171.460 116.045 171.630 ;
        RECT 111.200 171.130 111.370 171.320 ;
        RECT 116.340 171.130 116.510 171.320 ;
        RECT 111.665 170.820 116.045 170.990 ;
        RECT 111.200 170.490 111.370 170.680 ;
        RECT 116.340 170.490 116.510 170.680 ;
        RECT 111.665 170.180 116.045 170.350 ;
        RECT 111.200 169.850 111.370 170.040 ;
        RECT 116.340 169.850 116.510 170.040 ;
        RECT 111.665 169.540 116.045 169.710 ;
        RECT 111.200 169.210 111.370 169.400 ;
        RECT 116.340 169.210 116.510 169.400 ;
        RECT 111.665 168.900 116.045 169.070 ;
        RECT 111.200 168.570 111.370 168.760 ;
        RECT 116.340 168.570 116.510 168.760 ;
        RECT 111.665 168.260 116.045 168.430 ;
        RECT 111.200 167.930 111.370 168.120 ;
        RECT 116.340 167.930 116.510 168.120 ;
        RECT 111.665 167.620 116.045 167.790 ;
        RECT 111.200 167.290 111.370 167.480 ;
        RECT 116.340 167.290 116.510 167.480 ;
        RECT 111.665 166.980 116.045 167.150 ;
        RECT 111.200 166.650 111.370 166.840 ;
        RECT 116.340 166.650 116.510 166.840 ;
        RECT 111.665 166.340 116.045 166.510 ;
        RECT 111.200 166.010 111.370 166.200 ;
        RECT 116.340 166.010 116.510 166.200 ;
        RECT 111.665 165.700 116.045 165.870 ;
        RECT 111.200 165.370 111.370 165.560 ;
        RECT 116.340 165.370 116.510 165.560 ;
        RECT 111.665 165.060 116.045 165.230 ;
        RECT 111.200 164.730 111.370 164.920 ;
        RECT 116.340 164.730 116.510 164.920 ;
        RECT 111.665 164.420 116.045 164.590 ;
        RECT 111.200 164.090 111.370 164.280 ;
        RECT 116.340 164.090 116.510 164.280 ;
        RECT 111.665 163.780 116.045 163.950 ;
        RECT 111.200 163.450 111.370 163.640 ;
        RECT 116.340 163.450 116.510 163.640 ;
        RECT 111.665 163.140 116.045 163.310 ;
        RECT 111.200 162.810 111.370 163.000 ;
        RECT 116.340 162.810 116.510 163.000 ;
        RECT 111.665 162.500 116.045 162.670 ;
        RECT 111.200 162.170 111.370 162.360 ;
        RECT 116.340 162.170 116.510 162.360 ;
        RECT 111.665 161.860 116.045 162.030 ;
        RECT 111.200 161.530 111.370 161.720 ;
        RECT 116.340 161.530 116.510 161.720 ;
        RECT 111.665 161.220 116.045 161.390 ;
        RECT 111.200 160.890 111.370 161.080 ;
        RECT 116.340 160.890 116.510 161.080 ;
        RECT 111.665 160.580 116.045 160.750 ;
        RECT 111.200 160.250 111.370 160.440 ;
        RECT 116.340 160.250 116.510 160.440 ;
        RECT 111.665 159.940 116.045 160.110 ;
        RECT 111.200 159.610 111.370 159.800 ;
        RECT 116.340 159.610 116.510 159.800 ;
        RECT 111.665 159.300 116.045 159.470 ;
        RECT 111.200 158.970 111.370 159.160 ;
        RECT 116.340 158.970 116.510 159.160 ;
        RECT 111.665 158.660 116.045 158.830 ;
        RECT 117.320 157.730 117.490 173.430 ;
        RECT 118.250 157.730 118.420 173.430 ;
        RECT 119.635 173.040 121.015 173.210 ;
        RECT 119.170 172.800 119.340 172.970 ;
        RECT 121.310 172.800 121.480 172.970 ;
        RECT 119.635 172.560 121.015 172.730 ;
        RECT 119.170 172.320 119.340 172.490 ;
        RECT 121.310 172.320 121.480 172.490 ;
        RECT 119.635 172.080 121.015 172.250 ;
        RECT 130.520 173.570 131.210 173.740 ;
        RECT 119.635 170.940 121.015 171.110 ;
        RECT 119.170 170.700 119.340 170.870 ;
        RECT 121.310 170.700 121.480 170.870 ;
        RECT 119.635 170.460 121.015 170.630 ;
        RECT 119.170 170.220 119.340 170.390 ;
        RECT 121.310 170.220 121.480 170.390 ;
        RECT 119.635 169.980 121.015 170.150 ;
        RECT 123.480 172.520 124.860 172.690 ;
        RECT 123.060 172.300 123.230 172.470 ;
        RECT 125.110 172.300 125.280 172.470 ;
        RECT 123.480 172.080 124.860 172.250 ;
        RECT 126.170 172.430 127.170 173.430 ;
        RECT 123.480 170.940 124.860 171.110 ;
        RECT 123.060 170.720 123.230 170.890 ;
        RECT 125.110 170.720 125.280 170.890 ;
        RECT 123.480 170.500 124.860 170.670 ;
        RECT 120.080 167.080 124.460 167.250 ;
        RECT 119.660 166.750 119.830 166.940 ;
        RECT 124.710 166.750 124.880 166.940 ;
        RECT 120.080 166.440 124.460 166.610 ;
        RECT 119.660 166.110 119.830 166.300 ;
        RECT 124.710 166.110 124.880 166.300 ;
        RECT 120.080 165.800 124.460 165.970 ;
        RECT 119.660 165.470 119.830 165.660 ;
        RECT 124.710 165.470 124.880 165.660 ;
        RECT 120.080 165.160 124.460 165.330 ;
        RECT 119.660 164.830 119.830 165.020 ;
        RECT 124.710 164.830 124.880 165.020 ;
        RECT 120.080 164.520 124.460 164.690 ;
        RECT 119.660 164.190 119.830 164.380 ;
        RECT 124.710 164.190 124.880 164.380 ;
        RECT 120.080 163.880 124.460 164.050 ;
        RECT 119.660 163.550 119.830 163.740 ;
        RECT 124.710 163.550 124.880 163.740 ;
        RECT 120.080 163.240 124.460 163.410 ;
        RECT 119.660 162.910 119.830 163.100 ;
        RECT 124.710 162.910 124.880 163.100 ;
        RECT 120.080 162.600 124.460 162.770 ;
        RECT 117.370 156.430 118.370 157.430 ;
        RECT 126.120 156.430 126.290 172.130 ;
        RECT 130.770 171.005 130.960 172.990 ;
        RECT 130.770 158.850 130.960 160.835 ;
        RECT 134.765 172.210 139.145 172.380 ;
        RECT 134.300 171.880 134.470 172.070 ;
        RECT 139.440 171.880 139.610 172.070 ;
        RECT 134.765 171.570 139.145 171.740 ;
        RECT 134.300 171.240 134.470 171.430 ;
        RECT 139.440 171.240 139.610 171.430 ;
        RECT 134.765 170.930 139.145 171.100 ;
        RECT 134.300 170.600 134.470 170.790 ;
        RECT 139.440 170.600 139.610 170.790 ;
        RECT 134.765 170.290 139.145 170.460 ;
        RECT 134.300 169.960 134.470 170.150 ;
        RECT 139.440 169.960 139.610 170.150 ;
        RECT 134.765 169.650 139.145 169.820 ;
        RECT 134.300 169.320 134.470 169.510 ;
        RECT 139.440 169.320 139.610 169.510 ;
        RECT 134.765 169.010 139.145 169.180 ;
        RECT 134.300 168.680 134.470 168.870 ;
        RECT 139.440 168.680 139.610 168.870 ;
        RECT 134.765 168.370 139.145 168.540 ;
        RECT 134.300 168.040 134.470 168.230 ;
        RECT 139.440 168.040 139.610 168.230 ;
        RECT 134.765 167.730 139.145 167.900 ;
        RECT 134.300 167.400 134.470 167.590 ;
        RECT 139.440 167.400 139.610 167.590 ;
        RECT 134.765 167.090 139.145 167.260 ;
        RECT 134.300 166.760 134.470 166.950 ;
        RECT 139.440 166.760 139.610 166.950 ;
        RECT 134.765 166.450 139.145 166.620 ;
        RECT 134.300 166.120 134.470 166.310 ;
        RECT 139.440 166.120 139.610 166.310 ;
        RECT 134.765 165.810 139.145 165.980 ;
        RECT 134.300 165.480 134.470 165.670 ;
        RECT 139.440 165.480 139.610 165.670 ;
        RECT 134.765 165.170 139.145 165.340 ;
        RECT 134.300 164.840 134.470 165.030 ;
        RECT 139.440 164.840 139.610 165.030 ;
        RECT 134.765 164.530 139.145 164.700 ;
        RECT 134.300 164.200 134.470 164.390 ;
        RECT 139.440 164.200 139.610 164.390 ;
        RECT 134.765 163.890 139.145 164.060 ;
        RECT 134.300 163.560 134.470 163.750 ;
        RECT 139.440 163.560 139.610 163.750 ;
        RECT 134.765 163.250 139.145 163.420 ;
        RECT 134.300 162.920 134.470 163.110 ;
        RECT 139.440 162.920 139.610 163.110 ;
        RECT 134.765 162.610 139.145 162.780 ;
        RECT 134.300 162.280 134.470 162.470 ;
        RECT 139.440 162.280 139.610 162.470 ;
        RECT 134.765 161.970 139.145 162.140 ;
        RECT 134.300 161.640 134.470 161.830 ;
        RECT 139.440 161.640 139.610 161.830 ;
        RECT 134.765 161.330 139.145 161.500 ;
        RECT 134.300 161.000 134.470 161.190 ;
        RECT 139.440 161.000 139.610 161.190 ;
        RECT 134.765 160.690 139.145 160.860 ;
        RECT 134.300 160.360 134.470 160.550 ;
        RECT 139.440 160.360 139.610 160.550 ;
        RECT 134.765 160.050 139.145 160.220 ;
        RECT 134.300 159.720 134.470 159.910 ;
        RECT 139.440 159.720 139.610 159.910 ;
        RECT 134.765 159.410 139.145 159.580 ;
        RECT 134.300 159.080 134.470 159.270 ;
        RECT 139.440 159.080 139.610 159.270 ;
        RECT 134.765 158.770 139.145 158.940 ;
        RECT 140.420 157.840 140.590 173.540 ;
        RECT 141.350 157.840 141.520 173.540 ;
        RECT 142.735 173.150 144.115 173.320 ;
        RECT 142.270 172.910 142.440 173.080 ;
        RECT 144.410 172.910 144.580 173.080 ;
        RECT 142.735 172.670 144.115 172.840 ;
        RECT 142.270 172.430 142.440 172.600 ;
        RECT 144.410 172.430 144.580 172.600 ;
        RECT 142.735 172.190 144.115 172.360 ;
        RECT 142.735 171.050 144.115 171.220 ;
        RECT 142.270 170.810 142.440 170.980 ;
        RECT 144.410 170.810 144.580 170.980 ;
        RECT 142.735 170.570 144.115 170.740 ;
        RECT 142.270 170.330 142.440 170.500 ;
        RECT 144.410 170.330 144.580 170.500 ;
        RECT 142.735 170.090 144.115 170.260 ;
        RECT 146.580 172.630 147.960 172.800 ;
        RECT 146.160 172.410 146.330 172.580 ;
        RECT 148.210 172.410 148.380 172.580 ;
        RECT 146.580 172.190 147.960 172.360 ;
        RECT 149.270 172.540 150.270 173.540 ;
        RECT 146.580 171.050 147.960 171.220 ;
        RECT 146.160 170.830 146.330 171.000 ;
        RECT 148.210 170.830 148.380 171.000 ;
        RECT 146.580 170.610 147.960 170.780 ;
        RECT 143.180 167.190 147.560 167.360 ;
        RECT 142.760 166.860 142.930 167.050 ;
        RECT 147.810 166.860 147.980 167.050 ;
        RECT 143.180 166.550 147.560 166.720 ;
        RECT 142.760 166.220 142.930 166.410 ;
        RECT 147.810 166.220 147.980 166.410 ;
        RECT 143.180 165.910 147.560 166.080 ;
        RECT 142.760 165.580 142.930 165.770 ;
        RECT 147.810 165.580 147.980 165.770 ;
        RECT 143.180 165.270 147.560 165.440 ;
        RECT 142.760 164.940 142.930 165.130 ;
        RECT 147.810 164.940 147.980 165.130 ;
        RECT 143.180 164.630 147.560 164.800 ;
        RECT 142.760 164.300 142.930 164.490 ;
        RECT 147.810 164.300 147.980 164.490 ;
        RECT 143.180 163.990 147.560 164.160 ;
        RECT 142.760 163.660 142.930 163.850 ;
        RECT 147.810 163.660 147.980 163.850 ;
        RECT 143.180 163.350 147.560 163.520 ;
        RECT 142.760 163.020 142.930 163.210 ;
        RECT 147.810 163.020 147.980 163.210 ;
        RECT 143.180 162.710 147.560 162.880 ;
        RECT 140.470 156.540 141.470 157.540 ;
        RECT 149.220 156.540 149.390 172.240 ;
        RECT 84.730 147.620 85.420 147.790 ;
        RECT 84.980 145.055 85.170 147.040 ;
        RECT 84.980 132.900 85.170 134.885 ;
        RECT 88.975 146.260 93.355 146.430 ;
        RECT 88.510 145.930 88.680 146.120 ;
        RECT 93.650 145.930 93.820 146.120 ;
        RECT 88.975 145.620 93.355 145.790 ;
        RECT 88.510 145.290 88.680 145.480 ;
        RECT 93.650 145.290 93.820 145.480 ;
        RECT 88.975 144.980 93.355 145.150 ;
        RECT 88.510 144.650 88.680 144.840 ;
        RECT 93.650 144.650 93.820 144.840 ;
        RECT 88.975 144.340 93.355 144.510 ;
        RECT 88.510 144.010 88.680 144.200 ;
        RECT 93.650 144.010 93.820 144.200 ;
        RECT 88.975 143.700 93.355 143.870 ;
        RECT 88.510 143.370 88.680 143.560 ;
        RECT 93.650 143.370 93.820 143.560 ;
        RECT 88.975 143.060 93.355 143.230 ;
        RECT 88.510 142.730 88.680 142.920 ;
        RECT 93.650 142.730 93.820 142.920 ;
        RECT 88.975 142.420 93.355 142.590 ;
        RECT 88.510 142.090 88.680 142.280 ;
        RECT 93.650 142.090 93.820 142.280 ;
        RECT 88.975 141.780 93.355 141.950 ;
        RECT 88.510 141.450 88.680 141.640 ;
        RECT 93.650 141.450 93.820 141.640 ;
        RECT 88.975 141.140 93.355 141.310 ;
        RECT 88.510 140.810 88.680 141.000 ;
        RECT 93.650 140.810 93.820 141.000 ;
        RECT 88.975 140.500 93.355 140.670 ;
        RECT 88.510 140.170 88.680 140.360 ;
        RECT 93.650 140.170 93.820 140.360 ;
        RECT 88.975 139.860 93.355 140.030 ;
        RECT 88.510 139.530 88.680 139.720 ;
        RECT 93.650 139.530 93.820 139.720 ;
        RECT 88.975 139.220 93.355 139.390 ;
        RECT 88.510 138.890 88.680 139.080 ;
        RECT 93.650 138.890 93.820 139.080 ;
        RECT 88.975 138.580 93.355 138.750 ;
        RECT 88.510 138.250 88.680 138.440 ;
        RECT 93.650 138.250 93.820 138.440 ;
        RECT 88.975 137.940 93.355 138.110 ;
        RECT 88.510 137.610 88.680 137.800 ;
        RECT 93.650 137.610 93.820 137.800 ;
        RECT 88.975 137.300 93.355 137.470 ;
        RECT 88.510 136.970 88.680 137.160 ;
        RECT 93.650 136.970 93.820 137.160 ;
        RECT 88.975 136.660 93.355 136.830 ;
        RECT 88.510 136.330 88.680 136.520 ;
        RECT 93.650 136.330 93.820 136.520 ;
        RECT 88.975 136.020 93.355 136.190 ;
        RECT 88.510 135.690 88.680 135.880 ;
        RECT 93.650 135.690 93.820 135.880 ;
        RECT 88.975 135.380 93.355 135.550 ;
        RECT 88.510 135.050 88.680 135.240 ;
        RECT 93.650 135.050 93.820 135.240 ;
        RECT 88.975 134.740 93.355 134.910 ;
        RECT 88.510 134.410 88.680 134.600 ;
        RECT 93.650 134.410 93.820 134.600 ;
        RECT 88.975 134.100 93.355 134.270 ;
        RECT 88.510 133.770 88.680 133.960 ;
        RECT 93.650 133.770 93.820 133.960 ;
        RECT 88.975 133.460 93.355 133.630 ;
        RECT 88.510 133.130 88.680 133.320 ;
        RECT 93.650 133.130 93.820 133.320 ;
        RECT 88.975 132.820 93.355 132.990 ;
        RECT 94.630 131.890 94.800 147.590 ;
        RECT 95.560 131.890 95.730 147.590 ;
        RECT 96.945 147.200 98.325 147.370 ;
        RECT 96.480 146.960 96.650 147.130 ;
        RECT 98.620 146.960 98.790 147.130 ;
        RECT 96.945 146.720 98.325 146.890 ;
        RECT 96.480 146.480 96.650 146.650 ;
        RECT 98.620 146.480 98.790 146.650 ;
        RECT 96.945 146.240 98.325 146.410 ;
        RECT 107.760 147.770 108.450 147.940 ;
        RECT 96.945 145.100 98.325 145.270 ;
        RECT 96.480 144.860 96.650 145.030 ;
        RECT 98.620 144.860 98.790 145.030 ;
        RECT 96.945 144.620 98.325 144.790 ;
        RECT 96.480 144.380 96.650 144.550 ;
        RECT 98.620 144.380 98.790 144.550 ;
        RECT 96.945 144.140 98.325 144.310 ;
        RECT 100.790 146.680 102.170 146.850 ;
        RECT 100.370 146.460 100.540 146.630 ;
        RECT 102.420 146.460 102.590 146.630 ;
        RECT 100.790 146.240 102.170 146.410 ;
        RECT 103.480 146.590 104.480 147.590 ;
        RECT 100.790 145.100 102.170 145.270 ;
        RECT 100.370 144.880 100.540 145.050 ;
        RECT 102.420 144.880 102.590 145.050 ;
        RECT 100.790 144.660 102.170 144.830 ;
        RECT 97.390 141.240 101.770 141.410 ;
        RECT 96.970 140.910 97.140 141.100 ;
        RECT 102.020 140.910 102.190 141.100 ;
        RECT 97.390 140.600 101.770 140.770 ;
        RECT 96.970 140.270 97.140 140.460 ;
        RECT 102.020 140.270 102.190 140.460 ;
        RECT 97.390 139.960 101.770 140.130 ;
        RECT 96.970 139.630 97.140 139.820 ;
        RECT 102.020 139.630 102.190 139.820 ;
        RECT 97.390 139.320 101.770 139.490 ;
        RECT 96.970 138.990 97.140 139.180 ;
        RECT 102.020 138.990 102.190 139.180 ;
        RECT 97.390 138.680 101.770 138.850 ;
        RECT 96.970 138.350 97.140 138.540 ;
        RECT 102.020 138.350 102.190 138.540 ;
        RECT 97.390 138.040 101.770 138.210 ;
        RECT 96.970 137.710 97.140 137.900 ;
        RECT 102.020 137.710 102.190 137.900 ;
        RECT 97.390 137.400 101.770 137.570 ;
        RECT 96.970 137.070 97.140 137.260 ;
        RECT 102.020 137.070 102.190 137.260 ;
        RECT 97.390 136.760 101.770 136.930 ;
        RECT 94.680 130.590 95.680 131.590 ;
        RECT 103.430 130.590 103.600 146.290 ;
        RECT 108.010 145.205 108.200 147.190 ;
        RECT 108.010 133.050 108.200 135.035 ;
        RECT 112.005 146.410 116.385 146.580 ;
        RECT 111.540 146.080 111.710 146.270 ;
        RECT 116.680 146.080 116.850 146.270 ;
        RECT 112.005 145.770 116.385 145.940 ;
        RECT 111.540 145.440 111.710 145.630 ;
        RECT 116.680 145.440 116.850 145.630 ;
        RECT 112.005 145.130 116.385 145.300 ;
        RECT 111.540 144.800 111.710 144.990 ;
        RECT 116.680 144.800 116.850 144.990 ;
        RECT 112.005 144.490 116.385 144.660 ;
        RECT 111.540 144.160 111.710 144.350 ;
        RECT 116.680 144.160 116.850 144.350 ;
        RECT 112.005 143.850 116.385 144.020 ;
        RECT 111.540 143.520 111.710 143.710 ;
        RECT 116.680 143.520 116.850 143.710 ;
        RECT 112.005 143.210 116.385 143.380 ;
        RECT 111.540 142.880 111.710 143.070 ;
        RECT 116.680 142.880 116.850 143.070 ;
        RECT 112.005 142.570 116.385 142.740 ;
        RECT 111.540 142.240 111.710 142.430 ;
        RECT 116.680 142.240 116.850 142.430 ;
        RECT 112.005 141.930 116.385 142.100 ;
        RECT 111.540 141.600 111.710 141.790 ;
        RECT 116.680 141.600 116.850 141.790 ;
        RECT 112.005 141.290 116.385 141.460 ;
        RECT 111.540 140.960 111.710 141.150 ;
        RECT 116.680 140.960 116.850 141.150 ;
        RECT 112.005 140.650 116.385 140.820 ;
        RECT 111.540 140.320 111.710 140.510 ;
        RECT 116.680 140.320 116.850 140.510 ;
        RECT 112.005 140.010 116.385 140.180 ;
        RECT 111.540 139.680 111.710 139.870 ;
        RECT 116.680 139.680 116.850 139.870 ;
        RECT 112.005 139.370 116.385 139.540 ;
        RECT 111.540 139.040 111.710 139.230 ;
        RECT 116.680 139.040 116.850 139.230 ;
        RECT 112.005 138.730 116.385 138.900 ;
        RECT 111.540 138.400 111.710 138.590 ;
        RECT 116.680 138.400 116.850 138.590 ;
        RECT 112.005 138.090 116.385 138.260 ;
        RECT 111.540 137.760 111.710 137.950 ;
        RECT 116.680 137.760 116.850 137.950 ;
        RECT 112.005 137.450 116.385 137.620 ;
        RECT 111.540 137.120 111.710 137.310 ;
        RECT 116.680 137.120 116.850 137.310 ;
        RECT 112.005 136.810 116.385 136.980 ;
        RECT 111.540 136.480 111.710 136.670 ;
        RECT 116.680 136.480 116.850 136.670 ;
        RECT 112.005 136.170 116.385 136.340 ;
        RECT 111.540 135.840 111.710 136.030 ;
        RECT 116.680 135.840 116.850 136.030 ;
        RECT 112.005 135.530 116.385 135.700 ;
        RECT 111.540 135.200 111.710 135.390 ;
        RECT 116.680 135.200 116.850 135.390 ;
        RECT 112.005 134.890 116.385 135.060 ;
        RECT 111.540 134.560 111.710 134.750 ;
        RECT 116.680 134.560 116.850 134.750 ;
        RECT 112.005 134.250 116.385 134.420 ;
        RECT 111.540 133.920 111.710 134.110 ;
        RECT 116.680 133.920 116.850 134.110 ;
        RECT 112.005 133.610 116.385 133.780 ;
        RECT 111.540 133.280 111.710 133.470 ;
        RECT 116.680 133.280 116.850 133.470 ;
        RECT 112.005 132.970 116.385 133.140 ;
        RECT 117.660 132.040 117.830 147.740 ;
        RECT 118.590 132.040 118.760 147.740 ;
        RECT 119.975 147.350 121.355 147.520 ;
        RECT 119.510 147.110 119.680 147.280 ;
        RECT 121.650 147.110 121.820 147.280 ;
        RECT 119.975 146.870 121.355 147.040 ;
        RECT 119.510 146.630 119.680 146.800 ;
        RECT 121.650 146.630 121.820 146.800 ;
        RECT 119.975 146.390 121.355 146.560 ;
        RECT 130.770 147.850 131.460 148.020 ;
        RECT 119.975 145.250 121.355 145.420 ;
        RECT 119.510 145.010 119.680 145.180 ;
        RECT 121.650 145.010 121.820 145.180 ;
        RECT 119.975 144.770 121.355 144.940 ;
        RECT 119.510 144.530 119.680 144.700 ;
        RECT 121.650 144.530 121.820 144.700 ;
        RECT 119.975 144.290 121.355 144.460 ;
        RECT 123.820 146.830 125.200 147.000 ;
        RECT 123.400 146.610 123.570 146.780 ;
        RECT 125.450 146.610 125.620 146.780 ;
        RECT 123.820 146.390 125.200 146.560 ;
        RECT 126.510 146.740 127.510 147.740 ;
        RECT 123.820 145.250 125.200 145.420 ;
        RECT 123.400 145.030 123.570 145.200 ;
        RECT 125.450 145.030 125.620 145.200 ;
        RECT 123.820 144.810 125.200 144.980 ;
        RECT 120.420 141.390 124.800 141.560 ;
        RECT 120.000 141.060 120.170 141.250 ;
        RECT 125.050 141.060 125.220 141.250 ;
        RECT 120.420 140.750 124.800 140.920 ;
        RECT 120.000 140.420 120.170 140.610 ;
        RECT 125.050 140.420 125.220 140.610 ;
        RECT 120.420 140.110 124.800 140.280 ;
        RECT 120.000 139.780 120.170 139.970 ;
        RECT 125.050 139.780 125.220 139.970 ;
        RECT 120.420 139.470 124.800 139.640 ;
        RECT 120.000 139.140 120.170 139.330 ;
        RECT 125.050 139.140 125.220 139.330 ;
        RECT 120.420 138.830 124.800 139.000 ;
        RECT 120.000 138.500 120.170 138.690 ;
        RECT 125.050 138.500 125.220 138.690 ;
        RECT 120.420 138.190 124.800 138.360 ;
        RECT 120.000 137.860 120.170 138.050 ;
        RECT 125.050 137.860 125.220 138.050 ;
        RECT 120.420 137.550 124.800 137.720 ;
        RECT 120.000 137.220 120.170 137.410 ;
        RECT 125.050 137.220 125.220 137.410 ;
        RECT 120.420 136.910 124.800 137.080 ;
        RECT 117.710 130.740 118.710 131.740 ;
        RECT 126.460 130.740 126.630 146.440 ;
        RECT 131.020 145.285 131.210 147.270 ;
        RECT 131.020 133.130 131.210 135.115 ;
        RECT 135.015 146.490 139.395 146.660 ;
        RECT 134.550 146.160 134.720 146.350 ;
        RECT 139.690 146.160 139.860 146.350 ;
        RECT 135.015 145.850 139.395 146.020 ;
        RECT 134.550 145.520 134.720 145.710 ;
        RECT 139.690 145.520 139.860 145.710 ;
        RECT 135.015 145.210 139.395 145.380 ;
        RECT 134.550 144.880 134.720 145.070 ;
        RECT 139.690 144.880 139.860 145.070 ;
        RECT 135.015 144.570 139.395 144.740 ;
        RECT 134.550 144.240 134.720 144.430 ;
        RECT 139.690 144.240 139.860 144.430 ;
        RECT 135.015 143.930 139.395 144.100 ;
        RECT 134.550 143.600 134.720 143.790 ;
        RECT 139.690 143.600 139.860 143.790 ;
        RECT 135.015 143.290 139.395 143.460 ;
        RECT 134.550 142.960 134.720 143.150 ;
        RECT 139.690 142.960 139.860 143.150 ;
        RECT 135.015 142.650 139.395 142.820 ;
        RECT 134.550 142.320 134.720 142.510 ;
        RECT 139.690 142.320 139.860 142.510 ;
        RECT 135.015 142.010 139.395 142.180 ;
        RECT 134.550 141.680 134.720 141.870 ;
        RECT 139.690 141.680 139.860 141.870 ;
        RECT 135.015 141.370 139.395 141.540 ;
        RECT 134.550 141.040 134.720 141.230 ;
        RECT 139.690 141.040 139.860 141.230 ;
        RECT 135.015 140.730 139.395 140.900 ;
        RECT 134.550 140.400 134.720 140.590 ;
        RECT 139.690 140.400 139.860 140.590 ;
        RECT 135.015 140.090 139.395 140.260 ;
        RECT 134.550 139.760 134.720 139.950 ;
        RECT 139.690 139.760 139.860 139.950 ;
        RECT 135.015 139.450 139.395 139.620 ;
        RECT 134.550 139.120 134.720 139.310 ;
        RECT 139.690 139.120 139.860 139.310 ;
        RECT 135.015 138.810 139.395 138.980 ;
        RECT 134.550 138.480 134.720 138.670 ;
        RECT 139.690 138.480 139.860 138.670 ;
        RECT 135.015 138.170 139.395 138.340 ;
        RECT 134.550 137.840 134.720 138.030 ;
        RECT 139.690 137.840 139.860 138.030 ;
        RECT 135.015 137.530 139.395 137.700 ;
        RECT 134.550 137.200 134.720 137.390 ;
        RECT 139.690 137.200 139.860 137.390 ;
        RECT 135.015 136.890 139.395 137.060 ;
        RECT 134.550 136.560 134.720 136.750 ;
        RECT 139.690 136.560 139.860 136.750 ;
        RECT 135.015 136.250 139.395 136.420 ;
        RECT 134.550 135.920 134.720 136.110 ;
        RECT 139.690 135.920 139.860 136.110 ;
        RECT 135.015 135.610 139.395 135.780 ;
        RECT 134.550 135.280 134.720 135.470 ;
        RECT 139.690 135.280 139.860 135.470 ;
        RECT 135.015 134.970 139.395 135.140 ;
        RECT 134.550 134.640 134.720 134.830 ;
        RECT 139.690 134.640 139.860 134.830 ;
        RECT 135.015 134.330 139.395 134.500 ;
        RECT 134.550 134.000 134.720 134.190 ;
        RECT 139.690 134.000 139.860 134.190 ;
        RECT 135.015 133.690 139.395 133.860 ;
        RECT 134.550 133.360 134.720 133.550 ;
        RECT 139.690 133.360 139.860 133.550 ;
        RECT 135.015 133.050 139.395 133.220 ;
        RECT 140.670 132.120 140.840 147.820 ;
        RECT 141.600 132.120 141.770 147.820 ;
        RECT 142.985 147.430 144.365 147.600 ;
        RECT 142.520 147.190 142.690 147.360 ;
        RECT 144.660 147.190 144.830 147.360 ;
        RECT 142.985 146.950 144.365 147.120 ;
        RECT 142.520 146.710 142.690 146.880 ;
        RECT 144.660 146.710 144.830 146.880 ;
        RECT 142.985 146.470 144.365 146.640 ;
        RECT 142.985 145.330 144.365 145.500 ;
        RECT 142.520 145.090 142.690 145.260 ;
        RECT 144.660 145.090 144.830 145.260 ;
        RECT 142.985 144.850 144.365 145.020 ;
        RECT 142.520 144.610 142.690 144.780 ;
        RECT 144.660 144.610 144.830 144.780 ;
        RECT 142.985 144.370 144.365 144.540 ;
        RECT 146.830 146.910 148.210 147.080 ;
        RECT 146.410 146.690 146.580 146.860 ;
        RECT 148.460 146.690 148.630 146.860 ;
        RECT 146.830 146.470 148.210 146.640 ;
        RECT 149.520 146.820 150.520 147.820 ;
        RECT 146.830 145.330 148.210 145.500 ;
        RECT 146.410 145.110 146.580 145.280 ;
        RECT 148.460 145.110 148.630 145.280 ;
        RECT 146.830 144.890 148.210 145.060 ;
        RECT 143.430 141.470 147.810 141.640 ;
        RECT 143.010 141.140 143.180 141.330 ;
        RECT 148.060 141.140 148.230 141.330 ;
        RECT 143.430 140.830 147.810 141.000 ;
        RECT 143.010 140.500 143.180 140.690 ;
        RECT 148.060 140.500 148.230 140.690 ;
        RECT 143.430 140.190 147.810 140.360 ;
        RECT 143.010 139.860 143.180 140.050 ;
        RECT 148.060 139.860 148.230 140.050 ;
        RECT 143.430 139.550 147.810 139.720 ;
        RECT 143.010 139.220 143.180 139.410 ;
        RECT 148.060 139.220 148.230 139.410 ;
        RECT 143.430 138.910 147.810 139.080 ;
        RECT 143.010 138.580 143.180 138.770 ;
        RECT 148.060 138.580 148.230 138.770 ;
        RECT 143.430 138.270 147.810 138.440 ;
        RECT 143.010 137.940 143.180 138.130 ;
        RECT 148.060 137.940 148.230 138.130 ;
        RECT 143.430 137.630 147.810 137.800 ;
        RECT 143.010 137.300 143.180 137.490 ;
        RECT 148.060 137.300 148.230 137.490 ;
        RECT 143.430 136.990 147.810 137.160 ;
        RECT 140.720 130.820 141.720 131.820 ;
        RECT 149.470 130.820 149.640 146.520 ;
        RECT 58.610 34.050 59.450 34.220 ;
        RECT 57.740 24.020 57.910 33.310 ;
        RECT 58.300 23.875 58.470 33.755 ;
        RECT 59.590 23.875 59.760 33.755 ;
        RECT 58.610 23.410 59.450 23.580 ;
        RECT 58.560 16.570 59.400 16.740 ;
        RECT 57.680 6.630 57.850 16.050 ;
        RECT 58.250 6.440 58.420 16.320 ;
        RECT 59.540 6.440 59.710 16.320 ;
        RECT 58.560 6.020 59.400 6.190 ;
      LAYER met1 ;
        RECT 136.060 206.300 137.060 206.330 ;
        RECT 124.150 205.300 137.060 206.300 ;
        RECT 124.150 204.530 125.150 205.300 ;
        RECT 136.060 205.270 137.060 205.300 ;
        RECT 139.760 204.570 140.760 206.460 ;
        RECT 102.820 203.530 125.150 204.530 ;
        RECT 126.000 203.570 140.760 204.570 ;
        RECT 102.820 202.710 103.820 203.530 ;
        RECT 126.000 202.710 127.000 203.570 ;
        RECT 79.920 201.710 103.820 202.710 ;
        RECT 104.660 201.710 127.000 202.710 ;
        RECT 79.920 200.910 80.920 201.710 ;
        RECT 81.080 200.910 81.380 200.940 ;
        RECT 79.920 200.610 81.380 200.910 ;
        RECT 79.920 200.310 80.920 200.610 ;
        RECT 81.080 200.580 81.380 200.610 ;
        RECT 104.660 200.830 105.660 201.710 ;
        RECT 127.910 201.200 144.470 202.200 ;
        RECT 105.820 200.830 106.120 200.860 ;
        RECT 104.660 200.530 106.120 200.830 ;
        RECT 104.660 200.230 105.660 200.530 ;
        RECT 105.820 200.500 106.120 200.530 ;
        RECT 127.910 200.820 128.910 201.200 ;
        RECT 129.070 200.820 129.370 200.850 ;
        RECT 127.910 200.520 129.370 200.820 ;
        RECT 127.910 200.220 128.910 200.520 ;
        RECT 129.070 200.490 129.370 200.520 ;
        RECT 151.540 200.810 152.540 203.400 ;
        RECT 152.700 200.810 153.000 200.840 ;
        RECT 151.540 200.510 153.000 200.810 ;
        RECT 151.540 200.210 152.540 200.510 ;
        RECT 152.700 200.480 153.000 200.510 ;
        RECT 60.760 199.580 62.770 199.840 ;
        RECT 59.460 198.200 62.770 199.580 ;
        RECT 59.460 195.800 60.460 198.200 ;
        RECT 60.760 196.120 62.770 198.200 ;
        RECT 65.200 198.530 71.080 198.760 ;
        RECT 59.460 194.800 60.490 195.800 ;
        RECT 46.620 193.800 47.620 193.830 ;
        RECT 59.460 193.800 60.460 194.800 ;
        RECT 46.620 192.900 60.460 193.800 ;
        RECT 46.620 192.800 60.360 192.900 ;
        RECT 46.620 192.770 47.620 192.800 ;
        RECT 50.115 189.270 60.550 189.370 ;
        RECT 6.825 188.360 60.550 189.270 ;
        RECT 6.825 188.260 50.790 188.360 ;
        RECT 59.490 188.260 60.550 188.360 ;
        RECT 59.540 186.705 60.550 188.260 ;
        RECT 61.610 184.620 64.520 186.780 ;
        RECT 65.200 184.890 65.430 198.530 ;
        RECT 70.340 198.490 71.080 198.530 ;
        RECT 65.630 198.030 70.140 198.300 ;
        RECT 65.630 197.390 70.140 197.660 ;
        RECT 65.630 196.750 70.140 197.020 ;
        RECT 65.630 196.110 70.140 196.380 ;
        RECT 65.630 195.470 70.140 195.740 ;
        RECT 65.630 194.830 70.140 195.100 ;
        RECT 65.630 194.190 70.140 194.460 ;
        RECT 65.630 193.550 70.140 193.820 ;
        RECT 65.630 192.910 70.140 193.180 ;
        RECT 65.630 192.270 70.140 192.540 ;
        RECT 65.630 191.630 70.140 191.900 ;
        RECT 65.630 190.990 70.140 191.260 ;
        RECT 65.630 190.350 70.140 190.620 ;
        RECT 65.630 189.710 70.140 189.980 ;
        RECT 65.630 189.070 70.140 189.340 ;
        RECT 65.630 188.430 70.140 188.700 ;
        RECT 65.630 187.790 70.140 188.060 ;
        RECT 65.630 187.150 70.140 187.420 ;
        RECT 65.630 186.510 70.140 186.780 ;
        RECT 65.630 185.870 70.140 186.140 ;
        RECT 65.630 185.230 70.140 185.500 ;
        RECT 70.340 184.890 70.570 198.490 ;
        RECT 65.630 184.590 70.140 184.860 ;
        RECT 71.300 182.310 72.500 199.510 ;
        RECT 73.160 199.450 75.550 199.680 ;
        RECT 73.160 198.210 73.410 199.450 ;
        RECT 73.600 198.960 75.110 199.220 ;
        RECT 75.300 199.160 75.550 199.450 ;
        RECT 76.120 199.160 76.480 199.190 ;
        RECT 75.300 198.930 79.350 199.160 ;
        RECT 73.600 198.490 75.110 198.760 ;
        RECT 73.600 198.030 75.110 198.290 ;
        RECT 75.300 198.210 75.550 198.930 ;
        RECT 76.120 198.900 76.480 198.930 ;
        RECT 77.050 198.220 77.300 198.930 ;
        RECT 77.450 198.440 78.950 198.700 ;
        RECT 77.450 198.030 78.950 198.290 ;
        RECT 79.100 198.220 79.350 198.930 ;
        RECT 76.140 197.580 76.460 197.600 ;
        RECT 73.160 197.350 79.350 197.580 ;
        RECT 73.160 196.110 73.410 197.350 ;
        RECT 73.600 196.860 75.110 197.120 ;
        RECT 73.600 196.390 75.110 196.660 ;
        RECT 73.600 195.930 75.110 196.190 ;
        RECT 75.300 196.110 75.550 197.350 ;
        RECT 76.140 197.330 76.460 197.350 ;
        RECT 77.050 196.640 77.300 197.350 ;
        RECT 77.450 196.860 78.950 197.120 ;
        RECT 77.450 196.450 78.950 196.710 ;
        RECT 79.100 196.640 79.350 197.350 ;
        RECT 76.140 193.740 76.460 193.760 ;
        RECT 73.660 193.510 78.940 193.740 ;
        RECT 73.660 188.830 73.890 193.510 ;
        RECT 76.140 193.490 76.460 193.510 ;
        RECT 74.050 193.010 78.550 193.280 ;
        RECT 74.050 192.370 78.550 192.640 ;
        RECT 74.050 191.730 78.550 192.000 ;
        RECT 74.050 191.090 78.550 191.360 ;
        RECT 74.050 190.450 78.550 190.720 ;
        RECT 74.050 189.810 78.550 190.080 ;
        RECT 74.050 189.170 78.550 189.440 ;
        RECT 78.710 188.830 78.940 193.510 ;
        RECT 74.050 188.530 78.550 188.800 ;
        RECT 80.100 182.310 81.300 199.510 ;
        RECT 85.500 199.500 87.510 199.760 ;
        RECT 84.200 198.120 87.510 199.500 ;
        RECT 84.200 195.100 85.200 198.120 ;
        RECT 85.500 196.040 87.510 198.120 ;
        RECT 89.940 198.450 95.820 198.680 ;
        RECT 84.080 194.100 85.200 195.100 ;
        RECT 84.200 192.820 85.200 194.100 ;
        RECT 84.280 189.270 85.290 189.290 ;
        RECT 84.080 188.260 85.290 189.270 ;
        RECT 84.280 186.625 85.290 188.260 ;
        RECT 86.350 184.540 89.260 186.700 ;
        RECT 89.940 184.810 90.170 198.450 ;
        RECT 95.080 198.410 95.820 198.450 ;
        RECT 90.370 197.950 94.880 198.220 ;
        RECT 90.370 197.310 94.880 197.580 ;
        RECT 90.370 196.670 94.880 196.940 ;
        RECT 90.370 196.030 94.880 196.300 ;
        RECT 90.370 195.390 94.880 195.660 ;
        RECT 90.370 194.750 94.880 195.020 ;
        RECT 90.370 194.110 94.880 194.380 ;
        RECT 90.370 193.470 94.880 193.740 ;
        RECT 90.370 192.830 94.880 193.100 ;
        RECT 90.370 192.190 94.880 192.460 ;
        RECT 90.370 191.550 94.880 191.820 ;
        RECT 90.370 190.910 94.880 191.180 ;
        RECT 90.370 190.270 94.880 190.540 ;
        RECT 90.370 189.630 94.880 189.900 ;
        RECT 90.370 188.990 94.880 189.260 ;
        RECT 90.370 188.350 94.880 188.620 ;
        RECT 90.370 187.710 94.880 187.980 ;
        RECT 90.370 187.070 94.880 187.340 ;
        RECT 90.370 186.430 94.880 186.700 ;
        RECT 90.370 185.790 94.880 186.060 ;
        RECT 90.370 185.150 94.880 185.420 ;
        RECT 95.080 184.810 95.310 198.410 ;
        RECT 90.370 184.510 94.880 184.780 ;
        RECT 96.040 182.230 97.240 199.430 ;
        RECT 97.900 199.370 100.290 199.600 ;
        RECT 108.750 199.490 110.760 199.750 ;
        RECT 97.900 198.130 98.150 199.370 ;
        RECT 98.340 198.880 99.850 199.140 ;
        RECT 100.040 199.080 100.290 199.370 ;
        RECT 100.860 199.080 101.220 199.110 ;
        RECT 100.040 198.850 104.090 199.080 ;
        RECT 98.340 198.410 99.850 198.680 ;
        RECT 98.340 197.950 99.850 198.210 ;
        RECT 100.040 198.130 100.290 198.850 ;
        RECT 100.860 198.820 101.220 198.850 ;
        RECT 101.790 198.140 102.040 198.850 ;
        RECT 102.190 198.360 103.690 198.620 ;
        RECT 102.190 197.950 103.690 198.210 ;
        RECT 103.840 198.140 104.090 198.850 ;
        RECT 100.880 197.500 101.200 197.520 ;
        RECT 97.900 197.270 104.090 197.500 ;
        RECT 97.900 196.030 98.150 197.270 ;
        RECT 98.340 196.780 99.850 197.040 ;
        RECT 98.340 196.310 99.850 196.580 ;
        RECT 98.340 195.850 99.850 196.110 ;
        RECT 100.040 196.030 100.290 197.270 ;
        RECT 100.880 197.250 101.200 197.270 ;
        RECT 101.790 196.560 102.040 197.270 ;
        RECT 102.190 196.780 103.690 197.040 ;
        RECT 102.190 196.370 103.690 196.630 ;
        RECT 103.840 196.560 104.090 197.270 ;
        RECT 100.880 193.660 101.200 193.680 ;
        RECT 98.400 193.430 103.680 193.660 ;
        RECT 98.400 188.750 98.630 193.430 ;
        RECT 100.880 193.410 101.200 193.430 ;
        RECT 98.790 192.930 103.290 193.200 ;
        RECT 98.790 192.290 103.290 192.560 ;
        RECT 98.790 191.650 103.290 191.920 ;
        RECT 98.790 191.010 103.290 191.280 ;
        RECT 98.790 190.370 103.290 190.640 ;
        RECT 98.790 189.730 103.290 190.000 ;
        RECT 98.790 189.090 103.290 189.360 ;
        RECT 103.450 188.750 103.680 193.430 ;
        RECT 98.790 188.450 103.290 188.720 ;
        RECT 104.840 182.230 106.040 199.430 ;
        RECT 107.450 198.110 110.760 199.490 ;
        RECT 107.450 193.800 108.450 198.110 ;
        RECT 108.750 196.030 110.760 198.110 ;
        RECT 113.190 198.440 119.070 198.670 ;
        RECT 107.220 192.810 108.450 193.800 ;
        RECT 107.220 192.800 108.340 192.810 ;
        RECT 107.530 189.270 108.540 189.280 ;
        RECT 107.220 188.260 108.540 189.270 ;
        RECT 107.530 186.615 108.540 188.260 ;
        RECT 109.600 184.530 112.510 186.690 ;
        RECT 113.190 184.800 113.420 198.440 ;
        RECT 118.330 198.400 119.070 198.440 ;
        RECT 113.620 197.940 118.130 198.210 ;
        RECT 113.620 197.300 118.130 197.570 ;
        RECT 113.620 196.660 118.130 196.930 ;
        RECT 113.620 196.020 118.130 196.290 ;
        RECT 113.620 195.380 118.130 195.650 ;
        RECT 113.620 194.740 118.130 195.010 ;
        RECT 113.620 194.100 118.130 194.370 ;
        RECT 113.620 193.460 118.130 193.730 ;
        RECT 113.620 192.820 118.130 193.090 ;
        RECT 113.620 192.180 118.130 192.450 ;
        RECT 113.620 191.540 118.130 191.810 ;
        RECT 113.620 190.900 118.130 191.170 ;
        RECT 113.620 190.260 118.130 190.530 ;
        RECT 113.620 189.620 118.130 189.890 ;
        RECT 113.620 188.980 118.130 189.250 ;
        RECT 113.620 188.340 118.130 188.610 ;
        RECT 113.620 187.700 118.130 187.970 ;
        RECT 113.620 187.060 118.130 187.330 ;
        RECT 113.620 186.420 118.130 186.690 ;
        RECT 113.620 185.780 118.130 186.050 ;
        RECT 113.620 185.140 118.130 185.410 ;
        RECT 118.330 184.800 118.560 198.400 ;
        RECT 113.620 184.500 118.130 184.770 ;
        RECT 119.290 182.220 120.490 199.420 ;
        RECT 121.150 199.360 123.540 199.590 ;
        RECT 132.380 199.480 134.390 199.740 ;
        RECT 121.150 198.120 121.400 199.360 ;
        RECT 121.590 198.870 123.100 199.130 ;
        RECT 123.290 199.070 123.540 199.360 ;
        RECT 124.110 199.070 124.470 199.100 ;
        RECT 123.290 198.840 127.340 199.070 ;
        RECT 121.590 198.400 123.100 198.670 ;
        RECT 121.590 197.940 123.100 198.200 ;
        RECT 123.290 198.120 123.540 198.840 ;
        RECT 124.110 198.810 124.470 198.840 ;
        RECT 125.040 198.130 125.290 198.840 ;
        RECT 125.440 198.350 126.940 198.610 ;
        RECT 125.440 197.940 126.940 198.200 ;
        RECT 127.090 198.130 127.340 198.840 ;
        RECT 124.130 197.490 124.450 197.510 ;
        RECT 121.150 197.260 127.340 197.490 ;
        RECT 121.150 196.020 121.400 197.260 ;
        RECT 121.590 196.770 123.100 197.030 ;
        RECT 121.590 196.300 123.100 196.570 ;
        RECT 121.590 195.840 123.100 196.100 ;
        RECT 123.290 196.020 123.540 197.260 ;
        RECT 124.130 197.240 124.450 197.260 ;
        RECT 125.040 196.550 125.290 197.260 ;
        RECT 125.440 196.770 126.940 197.030 ;
        RECT 125.440 196.360 126.940 196.620 ;
        RECT 127.090 196.550 127.340 197.260 ;
        RECT 124.130 193.650 124.450 193.670 ;
        RECT 121.650 193.420 126.930 193.650 ;
        RECT 121.650 188.740 121.880 193.420 ;
        RECT 124.130 193.400 124.450 193.420 ;
        RECT 122.040 192.920 126.540 193.190 ;
        RECT 122.040 192.280 126.540 192.550 ;
        RECT 122.040 191.640 126.540 191.910 ;
        RECT 122.040 191.000 126.540 191.270 ;
        RECT 122.040 190.360 126.540 190.630 ;
        RECT 122.040 189.720 126.540 189.990 ;
        RECT 122.040 189.080 126.540 189.350 ;
        RECT 126.700 188.740 126.930 193.420 ;
        RECT 122.040 188.440 126.540 188.710 ;
        RECT 128.090 182.220 129.290 199.420 ;
        RECT 131.080 198.100 134.390 199.480 ;
        RECT 131.080 193.800 132.080 198.100 ;
        RECT 132.380 196.020 134.390 198.100 ;
        RECT 136.820 198.430 142.700 198.660 ;
        RECT 130.630 192.800 132.080 193.800 ;
        RECT 130.630 188.260 132.170 189.270 ;
        RECT 131.160 186.605 132.170 188.260 ;
        RECT 133.230 184.520 136.140 186.680 ;
        RECT 136.820 184.790 137.050 198.430 ;
        RECT 141.960 198.390 142.700 198.430 ;
        RECT 137.250 197.930 141.760 198.200 ;
        RECT 137.250 197.290 141.760 197.560 ;
        RECT 137.250 196.650 141.760 196.920 ;
        RECT 137.250 196.010 141.760 196.280 ;
        RECT 137.250 195.370 141.760 195.640 ;
        RECT 137.250 194.730 141.760 195.000 ;
        RECT 137.250 194.090 141.760 194.360 ;
        RECT 137.250 193.450 141.760 193.720 ;
        RECT 137.250 192.810 141.760 193.080 ;
        RECT 137.250 192.170 141.760 192.440 ;
        RECT 137.250 191.530 141.760 191.800 ;
        RECT 137.250 190.890 141.760 191.160 ;
        RECT 137.250 190.250 141.760 190.520 ;
        RECT 137.250 189.610 141.760 189.880 ;
        RECT 137.250 188.970 141.760 189.240 ;
        RECT 137.250 188.330 141.760 188.600 ;
        RECT 137.250 187.690 141.760 187.960 ;
        RECT 137.250 187.050 141.760 187.320 ;
        RECT 137.250 186.410 141.760 186.680 ;
        RECT 137.250 185.770 141.760 186.040 ;
        RECT 137.250 185.130 141.760 185.400 ;
        RECT 141.960 184.790 142.190 198.390 ;
        RECT 137.250 184.490 141.760 184.760 ;
        RECT 142.920 182.210 144.120 199.410 ;
        RECT 144.780 199.350 147.170 199.580 ;
        RECT 144.780 198.110 145.030 199.350 ;
        RECT 145.220 198.860 146.730 199.120 ;
        RECT 146.920 199.060 147.170 199.350 ;
        RECT 147.740 199.060 148.100 199.090 ;
        RECT 146.920 198.830 150.970 199.060 ;
        RECT 145.220 198.390 146.730 198.660 ;
        RECT 145.220 197.930 146.730 198.190 ;
        RECT 146.920 198.110 147.170 198.830 ;
        RECT 147.740 198.800 148.100 198.830 ;
        RECT 148.670 198.120 148.920 198.830 ;
        RECT 149.070 198.340 150.570 198.600 ;
        RECT 149.070 197.930 150.570 198.190 ;
        RECT 150.720 198.120 150.970 198.830 ;
        RECT 147.760 197.480 148.080 197.500 ;
        RECT 144.780 197.250 150.970 197.480 ;
        RECT 144.780 196.010 145.030 197.250 ;
        RECT 145.220 196.760 146.730 197.020 ;
        RECT 145.220 196.290 146.730 196.560 ;
        RECT 145.220 195.830 146.730 196.090 ;
        RECT 146.920 196.010 147.170 197.250 ;
        RECT 147.760 197.230 148.080 197.250 ;
        RECT 148.670 196.540 148.920 197.250 ;
        RECT 149.070 196.760 150.570 197.020 ;
        RECT 149.070 196.350 150.570 196.610 ;
        RECT 150.720 196.540 150.970 197.250 ;
        RECT 147.760 193.640 148.080 193.660 ;
        RECT 145.280 193.410 150.560 193.640 ;
        RECT 145.280 188.730 145.510 193.410 ;
        RECT 147.760 193.390 148.080 193.410 ;
        RECT 145.670 192.910 150.170 193.180 ;
        RECT 145.670 192.270 150.170 192.540 ;
        RECT 145.670 191.630 150.170 191.900 ;
        RECT 145.670 190.990 150.170 191.260 ;
        RECT 145.670 190.350 150.170 190.620 ;
        RECT 145.670 189.710 150.170 189.980 ;
        RECT 145.670 189.070 150.170 189.340 ;
        RECT 150.330 188.730 150.560 193.410 ;
        RECT 145.670 188.430 150.170 188.700 ;
        RECT 151.720 182.210 152.920 199.410 ;
        RECT 71.320 181.590 72.320 181.620 ;
        RECT 71.320 181.540 100.920 181.590 ;
        RECT 71.320 181.520 123.840 181.540 ;
        RECT 71.320 180.620 152.890 181.520 ;
        RECT 71.750 180.590 152.890 180.620 ;
        RECT 96.060 180.540 152.890 180.590 ;
        RECT 96.490 180.510 98.520 180.540 ;
        RECT 119.310 180.530 152.890 180.540 ;
        RECT 119.420 180.520 152.890 180.530 ;
        RECT 119.740 180.500 121.770 180.520 ;
        RECT 143.370 180.490 145.400 180.520 ;
        RECT 79.810 174.820 80.810 175.220 ;
        RECT 80.970 174.820 81.270 174.850 ;
        RECT 79.810 174.520 81.270 174.820 ;
        RECT 79.810 174.220 80.810 174.520 ;
        RECT 80.970 174.490 81.270 174.520 ;
        RECT 102.990 174.730 103.990 175.130 ;
        RECT 125.890 174.930 126.890 175.330 ;
        RECT 148.990 175.040 149.990 175.440 ;
        RECT 150.150 175.040 150.450 175.070 ;
        RECT 127.050 174.930 127.350 174.960 ;
        RECT 104.150 174.730 104.450 174.760 ;
        RECT 102.990 174.430 104.450 174.730 ;
        RECT 102.990 174.130 103.990 174.430 ;
        RECT 104.150 174.400 104.450 174.430 ;
        RECT 125.890 174.630 127.350 174.930 ;
        RECT 125.890 174.330 126.890 174.630 ;
        RECT 127.050 174.600 127.350 174.630 ;
        RECT 148.990 174.740 150.450 175.040 ;
        RECT 148.990 174.440 149.990 174.740 ;
        RECT 150.150 174.710 150.450 174.740 ;
        RECT 60.650 173.490 62.660 173.750 ;
        RECT 59.350 172.110 62.660 173.490 ;
        RECT 59.350 168.030 60.350 172.110 ;
        RECT 60.650 170.030 62.660 172.110 ;
        RECT 65.090 172.440 70.970 172.670 ;
        RECT 46.960 167.030 60.350 168.030 ;
        RECT 59.350 166.810 60.350 167.030 ;
        RECT 8.175 163.280 60.435 163.455 ;
        RECT 8.175 162.445 60.440 163.280 ;
        RECT 59.430 160.615 60.440 162.445 ;
        RECT 61.500 158.530 64.410 160.690 ;
        RECT 65.090 158.800 65.320 172.440 ;
        RECT 70.230 172.400 70.970 172.440 ;
        RECT 65.520 171.940 70.030 172.210 ;
        RECT 65.520 171.300 70.030 171.570 ;
        RECT 65.520 170.660 70.030 170.930 ;
        RECT 65.520 170.020 70.030 170.290 ;
        RECT 65.520 169.380 70.030 169.650 ;
        RECT 65.520 168.740 70.030 169.010 ;
        RECT 65.520 168.100 70.030 168.370 ;
        RECT 65.520 167.460 70.030 167.730 ;
        RECT 65.520 166.820 70.030 167.090 ;
        RECT 65.520 166.180 70.030 166.450 ;
        RECT 65.520 165.540 70.030 165.810 ;
        RECT 65.520 164.900 70.030 165.170 ;
        RECT 65.520 164.260 70.030 164.530 ;
        RECT 65.520 163.620 70.030 163.890 ;
        RECT 65.520 162.980 70.030 163.250 ;
        RECT 65.520 162.340 70.030 162.610 ;
        RECT 65.520 161.700 70.030 161.970 ;
        RECT 65.520 161.060 70.030 161.330 ;
        RECT 65.520 160.420 70.030 160.690 ;
        RECT 65.520 159.780 70.030 160.050 ;
        RECT 65.520 159.140 70.030 159.410 ;
        RECT 70.230 158.800 70.460 172.400 ;
        RECT 65.520 158.500 70.030 158.770 ;
        RECT 71.190 156.220 72.390 173.420 ;
        RECT 73.050 173.360 75.440 173.590 ;
        RECT 73.050 172.120 73.300 173.360 ;
        RECT 73.490 172.870 75.000 173.130 ;
        RECT 75.190 173.070 75.440 173.360 ;
        RECT 76.010 173.070 76.370 173.100 ;
        RECT 75.190 172.840 79.240 173.070 ;
        RECT 73.490 172.400 75.000 172.670 ;
        RECT 73.490 171.940 75.000 172.200 ;
        RECT 75.190 172.120 75.440 172.840 ;
        RECT 76.010 172.810 76.370 172.840 ;
        RECT 76.940 172.130 77.190 172.840 ;
        RECT 77.340 172.350 78.840 172.610 ;
        RECT 77.340 171.940 78.840 172.200 ;
        RECT 78.990 172.130 79.240 172.840 ;
        RECT 76.030 171.490 76.350 171.510 ;
        RECT 73.050 171.260 79.240 171.490 ;
        RECT 73.050 170.020 73.300 171.260 ;
        RECT 73.490 170.770 75.000 171.030 ;
        RECT 73.490 170.300 75.000 170.570 ;
        RECT 73.490 169.840 75.000 170.100 ;
        RECT 75.190 170.020 75.440 171.260 ;
        RECT 76.030 171.240 76.350 171.260 ;
        RECT 76.940 170.550 77.190 171.260 ;
        RECT 77.340 170.770 78.840 171.030 ;
        RECT 77.340 170.360 78.840 170.620 ;
        RECT 78.990 170.550 79.240 171.260 ;
        RECT 76.030 167.650 76.350 167.670 ;
        RECT 73.550 167.420 78.830 167.650 ;
        RECT 73.550 162.740 73.780 167.420 ;
        RECT 76.030 167.400 76.350 167.420 ;
        RECT 73.940 166.920 78.440 167.190 ;
        RECT 73.940 166.280 78.440 166.550 ;
        RECT 73.940 165.640 78.440 165.910 ;
        RECT 73.940 165.000 78.440 165.270 ;
        RECT 73.940 164.360 78.440 164.630 ;
        RECT 73.940 163.720 78.440 163.990 ;
        RECT 73.940 163.080 78.440 163.350 ;
        RECT 78.600 162.740 78.830 167.420 ;
        RECT 73.940 162.440 78.440 162.710 ;
        RECT 79.990 156.220 81.190 173.420 ;
        RECT 83.830 173.400 85.840 173.660 ;
        RECT 106.730 173.600 108.740 173.860 ;
        RECT 129.830 173.710 131.840 173.970 ;
        RECT 82.530 172.020 85.840 173.400 ;
        RECT 82.530 166.720 83.530 172.020 ;
        RECT 83.830 169.940 85.840 172.020 ;
        RECT 88.270 172.350 94.150 172.580 ;
        RECT 82.610 160.525 83.620 163.190 ;
        RECT 84.680 158.440 87.590 160.600 ;
        RECT 88.270 158.710 88.500 172.350 ;
        RECT 93.410 172.310 94.150 172.350 ;
        RECT 88.700 171.850 93.210 172.120 ;
        RECT 88.700 171.210 93.210 171.480 ;
        RECT 88.700 170.570 93.210 170.840 ;
        RECT 88.700 169.930 93.210 170.200 ;
        RECT 88.700 169.290 93.210 169.560 ;
        RECT 88.700 168.650 93.210 168.920 ;
        RECT 88.700 168.010 93.210 168.280 ;
        RECT 88.700 167.370 93.210 167.640 ;
        RECT 88.700 166.730 93.210 167.000 ;
        RECT 88.700 166.090 93.210 166.360 ;
        RECT 88.700 165.450 93.210 165.720 ;
        RECT 88.700 164.810 93.210 165.080 ;
        RECT 88.700 164.170 93.210 164.440 ;
        RECT 88.700 163.530 93.210 163.800 ;
        RECT 88.700 162.890 93.210 163.160 ;
        RECT 88.700 162.250 93.210 162.520 ;
        RECT 88.700 161.610 93.210 161.880 ;
        RECT 88.700 160.970 93.210 161.240 ;
        RECT 88.700 160.330 93.210 160.600 ;
        RECT 88.700 159.690 93.210 159.960 ;
        RECT 88.700 159.050 93.210 159.320 ;
        RECT 93.410 158.710 93.640 172.310 ;
        RECT 88.700 158.410 93.210 158.680 ;
        RECT 94.370 156.130 95.570 173.330 ;
        RECT 96.230 173.270 98.620 173.500 ;
        RECT 96.230 172.030 96.480 173.270 ;
        RECT 96.670 172.780 98.180 173.040 ;
        RECT 98.370 172.980 98.620 173.270 ;
        RECT 99.190 172.980 99.550 173.010 ;
        RECT 98.370 172.750 102.420 172.980 ;
        RECT 96.670 172.310 98.180 172.580 ;
        RECT 96.670 171.850 98.180 172.110 ;
        RECT 98.370 172.030 98.620 172.750 ;
        RECT 99.190 172.720 99.550 172.750 ;
        RECT 100.120 172.040 100.370 172.750 ;
        RECT 100.520 172.260 102.020 172.520 ;
        RECT 100.520 171.850 102.020 172.110 ;
        RECT 102.170 172.040 102.420 172.750 ;
        RECT 99.210 171.400 99.530 171.420 ;
        RECT 96.230 171.170 102.420 171.400 ;
        RECT 96.230 169.930 96.480 171.170 ;
        RECT 96.670 170.680 98.180 170.940 ;
        RECT 96.670 170.210 98.180 170.480 ;
        RECT 96.670 169.750 98.180 170.010 ;
        RECT 98.370 169.930 98.620 171.170 ;
        RECT 99.210 171.150 99.530 171.170 ;
        RECT 100.120 170.460 100.370 171.170 ;
        RECT 100.520 170.680 102.020 170.940 ;
        RECT 100.520 170.270 102.020 170.530 ;
        RECT 102.170 170.460 102.420 171.170 ;
        RECT 99.210 167.560 99.530 167.580 ;
        RECT 96.730 167.330 102.010 167.560 ;
        RECT 96.730 162.650 96.960 167.330 ;
        RECT 99.210 167.310 99.530 167.330 ;
        RECT 97.120 166.830 101.620 167.100 ;
        RECT 97.120 166.190 101.620 166.460 ;
        RECT 97.120 165.550 101.620 165.820 ;
        RECT 97.120 164.910 101.620 165.180 ;
        RECT 97.120 164.270 101.620 164.540 ;
        RECT 97.120 163.630 101.620 163.900 ;
        RECT 97.120 162.990 101.620 163.260 ;
        RECT 101.780 162.650 102.010 167.330 ;
        RECT 97.120 162.350 101.620 162.620 ;
        RECT 103.170 156.130 104.370 173.330 ;
        RECT 105.430 172.220 108.740 173.600 ;
        RECT 105.430 166.920 106.430 172.220 ;
        RECT 106.730 170.140 108.740 172.220 ;
        RECT 111.170 172.550 117.050 172.780 ;
        RECT 105.510 160.725 106.520 163.390 ;
        RECT 107.580 158.640 110.490 160.800 ;
        RECT 111.170 158.910 111.400 172.550 ;
        RECT 116.310 172.510 117.050 172.550 ;
        RECT 111.600 172.050 116.110 172.320 ;
        RECT 111.600 171.410 116.110 171.680 ;
        RECT 111.600 170.770 116.110 171.040 ;
        RECT 111.600 170.130 116.110 170.400 ;
        RECT 111.600 169.490 116.110 169.760 ;
        RECT 111.600 168.850 116.110 169.120 ;
        RECT 111.600 168.210 116.110 168.480 ;
        RECT 111.600 167.570 116.110 167.840 ;
        RECT 111.600 166.930 116.110 167.200 ;
        RECT 111.600 166.290 116.110 166.560 ;
        RECT 111.600 165.650 116.110 165.920 ;
        RECT 111.600 165.010 116.110 165.280 ;
        RECT 111.600 164.370 116.110 164.640 ;
        RECT 111.600 163.730 116.110 164.000 ;
        RECT 111.600 163.090 116.110 163.360 ;
        RECT 111.600 162.450 116.110 162.720 ;
        RECT 111.600 161.810 116.110 162.080 ;
        RECT 111.600 161.170 116.110 161.440 ;
        RECT 111.600 160.530 116.110 160.800 ;
        RECT 111.600 159.890 116.110 160.160 ;
        RECT 111.600 159.250 116.110 159.520 ;
        RECT 116.310 158.910 116.540 172.510 ;
        RECT 111.600 158.610 116.110 158.880 ;
        RECT 117.270 156.330 118.470 173.530 ;
        RECT 119.130 173.470 121.520 173.700 ;
        RECT 119.130 172.230 119.380 173.470 ;
        RECT 119.570 172.980 121.080 173.240 ;
        RECT 121.270 173.180 121.520 173.470 ;
        RECT 122.090 173.180 122.450 173.210 ;
        RECT 121.270 172.950 125.320 173.180 ;
        RECT 119.570 172.510 121.080 172.780 ;
        RECT 119.570 172.050 121.080 172.310 ;
        RECT 121.270 172.230 121.520 172.950 ;
        RECT 122.090 172.920 122.450 172.950 ;
        RECT 123.020 172.240 123.270 172.950 ;
        RECT 123.420 172.460 124.920 172.720 ;
        RECT 123.420 172.050 124.920 172.310 ;
        RECT 125.070 172.240 125.320 172.950 ;
        RECT 122.110 171.600 122.430 171.620 ;
        RECT 119.130 171.370 125.320 171.600 ;
        RECT 119.130 170.130 119.380 171.370 ;
        RECT 119.570 170.880 121.080 171.140 ;
        RECT 119.570 170.410 121.080 170.680 ;
        RECT 119.570 169.950 121.080 170.210 ;
        RECT 121.270 170.130 121.520 171.370 ;
        RECT 122.110 171.350 122.430 171.370 ;
        RECT 123.020 170.660 123.270 171.370 ;
        RECT 123.420 170.880 124.920 171.140 ;
        RECT 123.420 170.470 124.920 170.730 ;
        RECT 125.070 170.660 125.320 171.370 ;
        RECT 122.110 167.760 122.430 167.780 ;
        RECT 119.630 167.530 124.910 167.760 ;
        RECT 119.630 162.850 119.860 167.530 ;
        RECT 122.110 167.510 122.430 167.530 ;
        RECT 120.020 167.030 124.520 167.300 ;
        RECT 120.020 166.390 124.520 166.660 ;
        RECT 120.020 165.750 124.520 166.020 ;
        RECT 120.020 165.110 124.520 165.380 ;
        RECT 120.020 164.470 124.520 164.740 ;
        RECT 120.020 163.830 124.520 164.100 ;
        RECT 120.020 163.190 124.520 163.460 ;
        RECT 124.680 162.850 124.910 167.530 ;
        RECT 120.020 162.550 124.520 162.820 ;
        RECT 126.070 156.330 127.270 173.530 ;
        RECT 128.530 172.330 131.840 173.710 ;
        RECT 128.530 167.030 129.530 172.330 ;
        RECT 129.830 170.250 131.840 172.330 ;
        RECT 134.270 172.660 140.150 172.890 ;
        RECT 128.610 160.835 129.620 163.500 ;
        RECT 130.680 158.750 133.590 160.910 ;
        RECT 134.270 159.020 134.500 172.660 ;
        RECT 139.410 172.620 140.150 172.660 ;
        RECT 134.700 172.160 139.210 172.430 ;
        RECT 134.700 171.520 139.210 171.790 ;
        RECT 134.700 170.880 139.210 171.150 ;
        RECT 134.700 170.240 139.210 170.510 ;
        RECT 134.700 169.600 139.210 169.870 ;
        RECT 134.700 168.960 139.210 169.230 ;
        RECT 134.700 168.320 139.210 168.590 ;
        RECT 134.700 167.680 139.210 167.950 ;
        RECT 134.700 167.040 139.210 167.310 ;
        RECT 134.700 166.400 139.210 166.670 ;
        RECT 134.700 165.760 139.210 166.030 ;
        RECT 134.700 165.120 139.210 165.390 ;
        RECT 134.700 164.480 139.210 164.750 ;
        RECT 134.700 163.840 139.210 164.110 ;
        RECT 134.700 163.200 139.210 163.470 ;
        RECT 134.700 162.560 139.210 162.830 ;
        RECT 134.700 161.920 139.210 162.190 ;
        RECT 134.700 161.280 139.210 161.550 ;
        RECT 134.700 160.640 139.210 160.910 ;
        RECT 134.700 160.000 139.210 160.270 ;
        RECT 134.700 159.360 139.210 159.630 ;
        RECT 139.410 159.020 139.640 172.620 ;
        RECT 134.700 158.720 139.210 158.990 ;
        RECT 140.370 156.440 141.570 173.640 ;
        RECT 142.230 173.580 144.620 173.810 ;
        RECT 142.230 172.340 142.480 173.580 ;
        RECT 142.670 173.090 144.180 173.350 ;
        RECT 144.370 173.290 144.620 173.580 ;
        RECT 145.190 173.290 145.550 173.320 ;
        RECT 144.370 173.060 148.420 173.290 ;
        RECT 142.670 172.620 144.180 172.890 ;
        RECT 142.670 172.160 144.180 172.420 ;
        RECT 144.370 172.340 144.620 173.060 ;
        RECT 145.190 173.030 145.550 173.060 ;
        RECT 146.120 172.350 146.370 173.060 ;
        RECT 146.520 172.570 148.020 172.830 ;
        RECT 146.520 172.160 148.020 172.420 ;
        RECT 148.170 172.350 148.420 173.060 ;
        RECT 145.210 171.710 145.530 171.730 ;
        RECT 142.230 171.480 148.420 171.710 ;
        RECT 142.230 170.240 142.480 171.480 ;
        RECT 142.670 170.990 144.180 171.250 ;
        RECT 142.670 170.520 144.180 170.790 ;
        RECT 142.670 170.060 144.180 170.320 ;
        RECT 144.370 170.240 144.620 171.480 ;
        RECT 145.210 171.460 145.530 171.480 ;
        RECT 146.120 170.770 146.370 171.480 ;
        RECT 146.520 170.990 148.020 171.250 ;
        RECT 146.520 170.580 148.020 170.840 ;
        RECT 148.170 170.770 148.420 171.480 ;
        RECT 145.210 167.870 145.530 167.890 ;
        RECT 142.730 167.640 148.010 167.870 ;
        RECT 142.730 162.960 142.960 167.640 ;
        RECT 145.210 167.620 145.530 167.640 ;
        RECT 143.120 167.140 147.620 167.410 ;
        RECT 143.120 166.500 147.620 166.770 ;
        RECT 143.120 165.860 147.620 166.130 ;
        RECT 143.120 165.220 147.620 165.490 ;
        RECT 143.120 164.580 147.620 164.850 ;
        RECT 143.120 163.940 147.620 164.210 ;
        RECT 143.120 163.300 147.620 163.570 ;
        RECT 147.780 162.960 148.010 167.640 ;
        RECT 143.120 162.660 147.620 162.930 ;
        RECT 149.170 156.440 150.370 173.640 ;
        RECT 140.390 155.720 141.390 155.750 ;
        RECT 117.290 155.610 118.290 155.640 ;
        RECT 140.390 155.610 142.850 155.720 ;
        RECT 71.210 155.440 95.380 155.530 ;
        RECT 71.210 155.410 95.390 155.440 ;
        RECT 117.290 155.410 142.850 155.610 ;
        RECT 71.210 154.720 142.850 155.410 ;
        RECT 71.210 154.610 141.380 154.720 ;
        RECT 71.210 154.530 118.250 154.610 ;
        RECT 71.640 154.500 73.670 154.530 ;
        RECT 94.390 154.440 118.250 154.530 ;
        RECT 94.820 154.410 118.250 154.440 ;
        RECT 103.200 149.090 104.200 149.490 ;
        RECT 126.230 149.240 127.230 149.640 ;
        RECT 149.240 149.320 150.240 149.720 ;
        RECT 150.400 149.320 150.700 149.350 ;
        RECT 127.390 149.240 127.690 149.270 ;
        RECT 104.360 149.090 104.660 149.120 ;
        RECT 103.200 148.790 104.660 149.090 ;
        RECT 103.200 148.490 104.200 148.790 ;
        RECT 104.360 148.760 104.660 148.790 ;
        RECT 126.230 148.940 127.690 149.240 ;
        RECT 126.230 148.640 127.230 148.940 ;
        RECT 127.390 148.910 127.690 148.940 ;
        RECT 149.240 149.020 150.700 149.320 ;
        RECT 149.240 148.720 150.240 149.020 ;
        RECT 150.400 148.990 150.700 149.020 ;
        RECT 84.040 147.760 86.050 148.020 ;
        RECT 107.070 147.910 109.080 148.170 ;
        RECT 82.740 146.380 86.050 147.760 ;
        RECT 82.740 142.310 83.740 146.380 ;
        RECT 84.040 144.300 86.050 146.380 ;
        RECT 88.480 146.710 94.360 146.940 ;
        RECT 57.140 141.310 83.740 142.310 ;
        RECT 82.740 141.080 83.740 141.310 ;
        RECT 8.235 137.550 83.785 137.780 ;
        RECT 8.235 136.770 83.830 137.550 ;
        RECT 82.820 134.885 83.830 136.770 ;
        RECT 84.890 132.800 87.800 134.960 ;
        RECT 88.480 133.070 88.710 146.710 ;
        RECT 93.620 146.670 94.360 146.710 ;
        RECT 88.910 146.210 93.420 146.480 ;
        RECT 88.910 145.570 93.420 145.840 ;
        RECT 88.910 144.930 93.420 145.200 ;
        RECT 88.910 144.290 93.420 144.560 ;
        RECT 88.910 143.650 93.420 143.920 ;
        RECT 88.910 143.010 93.420 143.280 ;
        RECT 88.910 142.370 93.420 142.640 ;
        RECT 88.910 141.730 93.420 142.000 ;
        RECT 88.910 141.090 93.420 141.360 ;
        RECT 88.910 140.450 93.420 140.720 ;
        RECT 88.910 139.810 93.420 140.080 ;
        RECT 88.910 139.170 93.420 139.440 ;
        RECT 88.910 138.530 93.420 138.800 ;
        RECT 88.910 137.890 93.420 138.160 ;
        RECT 88.910 137.250 93.420 137.520 ;
        RECT 88.910 136.610 93.420 136.880 ;
        RECT 88.910 135.970 93.420 136.240 ;
        RECT 88.910 135.330 93.420 135.600 ;
        RECT 88.910 134.690 93.420 134.960 ;
        RECT 88.910 134.050 93.420 134.320 ;
        RECT 88.910 133.410 93.420 133.680 ;
        RECT 93.620 133.070 93.850 146.670 ;
        RECT 88.910 132.770 93.420 133.040 ;
        RECT 94.580 130.490 95.780 147.690 ;
        RECT 96.440 147.630 98.830 147.860 ;
        RECT 96.440 146.390 96.690 147.630 ;
        RECT 96.880 147.140 98.390 147.400 ;
        RECT 98.580 147.340 98.830 147.630 ;
        RECT 99.400 147.340 99.760 147.370 ;
        RECT 98.580 147.110 102.630 147.340 ;
        RECT 96.880 146.670 98.390 146.940 ;
        RECT 96.880 146.210 98.390 146.470 ;
        RECT 98.580 146.390 98.830 147.110 ;
        RECT 99.400 147.080 99.760 147.110 ;
        RECT 100.330 146.400 100.580 147.110 ;
        RECT 100.730 146.620 102.230 146.880 ;
        RECT 100.730 146.210 102.230 146.470 ;
        RECT 102.380 146.400 102.630 147.110 ;
        RECT 99.420 145.760 99.740 145.780 ;
        RECT 96.440 145.530 102.630 145.760 ;
        RECT 96.440 144.290 96.690 145.530 ;
        RECT 96.880 145.040 98.390 145.300 ;
        RECT 96.880 144.570 98.390 144.840 ;
        RECT 96.880 144.110 98.390 144.370 ;
        RECT 98.580 144.290 98.830 145.530 ;
        RECT 99.420 145.510 99.740 145.530 ;
        RECT 100.330 144.820 100.580 145.530 ;
        RECT 100.730 145.040 102.230 145.300 ;
        RECT 100.730 144.630 102.230 144.890 ;
        RECT 102.380 144.820 102.630 145.530 ;
        RECT 99.420 141.920 99.740 141.940 ;
        RECT 96.940 141.690 102.220 141.920 ;
        RECT 96.940 137.010 97.170 141.690 ;
        RECT 99.420 141.670 99.740 141.690 ;
        RECT 97.330 141.190 101.830 141.460 ;
        RECT 97.330 140.550 101.830 140.820 ;
        RECT 97.330 139.910 101.830 140.180 ;
        RECT 97.330 139.270 101.830 139.540 ;
        RECT 97.330 138.630 101.830 138.900 ;
        RECT 97.330 137.990 101.830 138.260 ;
        RECT 97.330 137.350 101.830 137.620 ;
        RECT 101.990 137.010 102.220 141.690 ;
        RECT 97.330 136.710 101.830 136.980 ;
        RECT 103.380 130.490 104.580 147.690 ;
        RECT 105.770 146.530 109.080 147.910 ;
        RECT 105.770 141.230 106.770 146.530 ;
        RECT 107.070 144.450 109.080 146.530 ;
        RECT 111.510 146.860 117.390 147.090 ;
        RECT 105.850 135.035 106.860 137.700 ;
        RECT 107.920 132.950 110.830 135.110 ;
        RECT 111.510 133.220 111.740 146.860 ;
        RECT 116.650 146.820 117.390 146.860 ;
        RECT 111.940 146.360 116.450 146.630 ;
        RECT 111.940 145.720 116.450 145.990 ;
        RECT 111.940 145.080 116.450 145.350 ;
        RECT 111.940 144.440 116.450 144.710 ;
        RECT 111.940 143.800 116.450 144.070 ;
        RECT 111.940 143.160 116.450 143.430 ;
        RECT 111.940 142.520 116.450 142.790 ;
        RECT 111.940 141.880 116.450 142.150 ;
        RECT 111.940 141.240 116.450 141.510 ;
        RECT 111.940 140.600 116.450 140.870 ;
        RECT 111.940 139.960 116.450 140.230 ;
        RECT 111.940 139.320 116.450 139.590 ;
        RECT 111.940 138.680 116.450 138.950 ;
        RECT 111.940 138.040 116.450 138.310 ;
        RECT 111.940 137.400 116.450 137.670 ;
        RECT 111.940 136.760 116.450 137.030 ;
        RECT 111.940 136.120 116.450 136.390 ;
        RECT 111.940 135.480 116.450 135.750 ;
        RECT 111.940 134.840 116.450 135.110 ;
        RECT 111.940 134.200 116.450 134.470 ;
        RECT 111.940 133.560 116.450 133.830 ;
        RECT 116.650 133.220 116.880 146.820 ;
        RECT 111.940 132.920 116.450 133.190 ;
        RECT 117.610 130.640 118.810 147.840 ;
        RECT 119.470 147.780 121.860 148.010 ;
        RECT 130.080 147.990 132.090 148.250 ;
        RECT 119.470 146.540 119.720 147.780 ;
        RECT 119.910 147.290 121.420 147.550 ;
        RECT 121.610 147.490 121.860 147.780 ;
        RECT 122.430 147.490 122.790 147.520 ;
        RECT 121.610 147.260 125.660 147.490 ;
        RECT 119.910 146.820 121.420 147.090 ;
        RECT 119.910 146.360 121.420 146.620 ;
        RECT 121.610 146.540 121.860 147.260 ;
        RECT 122.430 147.230 122.790 147.260 ;
        RECT 123.360 146.550 123.610 147.260 ;
        RECT 123.760 146.770 125.260 147.030 ;
        RECT 123.760 146.360 125.260 146.620 ;
        RECT 125.410 146.550 125.660 147.260 ;
        RECT 122.450 145.910 122.770 145.930 ;
        RECT 119.470 145.680 125.660 145.910 ;
        RECT 119.470 144.440 119.720 145.680 ;
        RECT 119.910 145.190 121.420 145.450 ;
        RECT 119.910 144.720 121.420 144.990 ;
        RECT 119.910 144.260 121.420 144.520 ;
        RECT 121.610 144.440 121.860 145.680 ;
        RECT 122.450 145.660 122.770 145.680 ;
        RECT 123.360 144.970 123.610 145.680 ;
        RECT 123.760 145.190 125.260 145.450 ;
        RECT 123.760 144.780 125.260 145.040 ;
        RECT 125.410 144.970 125.660 145.680 ;
        RECT 122.450 142.070 122.770 142.090 ;
        RECT 119.970 141.840 125.250 142.070 ;
        RECT 119.970 137.160 120.200 141.840 ;
        RECT 122.450 141.820 122.770 141.840 ;
        RECT 120.360 141.340 124.860 141.610 ;
        RECT 120.360 140.700 124.860 140.970 ;
        RECT 120.360 140.060 124.860 140.330 ;
        RECT 120.360 139.420 124.860 139.690 ;
        RECT 120.360 138.780 124.860 139.050 ;
        RECT 120.360 138.140 124.860 138.410 ;
        RECT 120.360 137.500 124.860 137.770 ;
        RECT 125.020 137.160 125.250 141.840 ;
        RECT 120.360 136.860 124.860 137.130 ;
        RECT 126.410 130.640 127.610 147.840 ;
        RECT 128.780 146.610 132.090 147.990 ;
        RECT 128.780 141.310 129.780 146.610 ;
        RECT 130.080 144.530 132.090 146.610 ;
        RECT 134.520 146.940 140.400 147.170 ;
        RECT 128.860 135.115 129.870 137.780 ;
        RECT 130.930 133.030 133.840 135.190 ;
        RECT 134.520 133.300 134.750 146.940 ;
        RECT 139.660 146.900 140.400 146.940 ;
        RECT 134.950 146.440 139.460 146.710 ;
        RECT 134.950 145.800 139.460 146.070 ;
        RECT 134.950 145.160 139.460 145.430 ;
        RECT 134.950 144.520 139.460 144.790 ;
        RECT 134.950 143.880 139.460 144.150 ;
        RECT 134.950 143.240 139.460 143.510 ;
        RECT 134.950 142.600 139.460 142.870 ;
        RECT 134.950 141.960 139.460 142.230 ;
        RECT 134.950 141.320 139.460 141.590 ;
        RECT 134.950 140.680 139.460 140.950 ;
        RECT 134.950 140.040 139.460 140.310 ;
        RECT 134.950 139.400 139.460 139.670 ;
        RECT 134.950 138.760 139.460 139.030 ;
        RECT 134.950 138.120 139.460 138.390 ;
        RECT 134.950 137.480 139.460 137.750 ;
        RECT 134.950 136.840 139.460 137.110 ;
        RECT 134.950 136.200 139.460 136.470 ;
        RECT 134.950 135.560 139.460 135.830 ;
        RECT 134.950 134.920 139.460 135.190 ;
        RECT 134.950 134.280 139.460 134.550 ;
        RECT 134.950 133.640 139.460 133.910 ;
        RECT 139.660 133.300 139.890 146.900 ;
        RECT 134.950 133.000 139.460 133.270 ;
        RECT 140.620 130.720 141.820 147.920 ;
        RECT 142.480 147.860 144.870 148.090 ;
        RECT 142.480 146.620 142.730 147.860 ;
        RECT 142.920 147.370 144.430 147.630 ;
        RECT 144.620 147.570 144.870 147.860 ;
        RECT 145.440 147.570 145.800 147.600 ;
        RECT 144.620 147.340 148.670 147.570 ;
        RECT 142.920 146.900 144.430 147.170 ;
        RECT 142.920 146.440 144.430 146.700 ;
        RECT 144.620 146.620 144.870 147.340 ;
        RECT 145.440 147.310 145.800 147.340 ;
        RECT 146.370 146.630 146.620 147.340 ;
        RECT 146.770 146.850 148.270 147.110 ;
        RECT 146.770 146.440 148.270 146.700 ;
        RECT 148.420 146.630 148.670 147.340 ;
        RECT 145.460 145.990 145.780 146.010 ;
        RECT 142.480 145.760 148.670 145.990 ;
        RECT 142.480 144.520 142.730 145.760 ;
        RECT 142.920 145.270 144.430 145.530 ;
        RECT 142.920 144.800 144.430 145.070 ;
        RECT 142.920 144.340 144.430 144.600 ;
        RECT 144.620 144.520 144.870 145.760 ;
        RECT 145.460 145.740 145.780 145.760 ;
        RECT 146.370 145.050 146.620 145.760 ;
        RECT 146.770 145.270 148.270 145.530 ;
        RECT 146.770 144.860 148.270 145.120 ;
        RECT 148.420 145.050 148.670 145.760 ;
        RECT 145.460 142.150 145.780 142.170 ;
        RECT 142.980 141.920 148.260 142.150 ;
        RECT 142.980 137.240 143.210 141.920 ;
        RECT 145.460 141.900 145.780 141.920 ;
        RECT 143.370 141.420 147.870 141.690 ;
        RECT 143.370 140.780 147.870 141.050 ;
        RECT 143.370 140.140 147.870 140.410 ;
        RECT 143.370 139.500 147.870 139.770 ;
        RECT 143.370 138.860 147.870 139.130 ;
        RECT 143.370 138.220 147.870 138.490 ;
        RECT 143.370 137.580 147.870 137.850 ;
        RECT 148.030 137.240 148.260 141.920 ;
        RECT 143.370 136.940 147.870 137.210 ;
        RECT 149.420 130.720 150.620 147.920 ;
        RECT 117.750 130.000 141.640 130.030 ;
        RECT 117.750 129.950 143.100 130.000 ;
        RECT 117.630 129.800 143.100 129.950 ;
        RECT 94.600 129.030 143.100 129.800 ;
        RECT 94.600 128.800 122.210 129.030 ;
        RECT 141.070 129.000 143.100 129.030 ;
        RECT 95.030 128.770 97.060 128.800 ;
        RECT 53.345 34.530 59.530 35.530 ;
        RECT 53.345 34.220 54.345 34.530 ;
        RECT 53.345 34.050 54.350 34.220 ;
        RECT 53.345 23.580 54.345 34.050 ;
        RECT 58.530 33.980 59.530 34.530 ;
        RECT 55.230 33.660 57.210 33.770 ;
        RECT 58.270 33.660 58.500 33.815 ;
        RECT 55.230 24.020 58.500 33.660 ;
        RECT 55.230 23.870 57.420 24.020 ;
        RECT 57.710 23.980 57.970 24.020 ;
        RECT 57.710 23.970 57.930 23.980 ;
        RECT 58.270 23.815 58.500 24.020 ;
        RECT 59.560 33.760 59.790 33.815 ;
        RECT 59.560 23.870 61.580 33.760 ;
        RECT 59.560 23.815 59.790 23.870 ;
        RECT 53.345 23.410 54.350 23.580 ;
        RECT 53.345 20.490 54.345 23.410 ;
        RECT 51.245 20.330 54.350 20.490 ;
        RECT 58.540 20.410 59.540 23.610 ;
        RECT 60.590 20.535 61.580 23.870 ;
        RECT 58.530 20.330 59.550 20.410 ;
        RECT 51.245 19.330 59.550 20.330 ;
        RECT 51.245 19.165 54.350 19.330 ;
        RECT 53.345 5.420 54.345 19.165 ;
        RECT 58.530 16.770 59.550 19.330 ;
        RECT 60.395 19.105 61.765 20.535 ;
        RECT 60.590 18.395 61.580 19.105 ;
        RECT 58.500 16.540 59.550 16.770 ;
        RECT 55.230 16.050 57.280 16.280 ;
        RECT 57.620 16.050 57.880 16.110 ;
        RECT 58.220 16.050 58.450 16.380 ;
        RECT 55.230 6.560 58.450 16.050 ;
        RECT 55.230 6.480 57.340 6.560 ;
        RECT 55.230 6.460 57.300 6.480 ;
        RECT 58.220 6.380 58.450 6.560 ;
        RECT 59.510 16.280 59.740 16.380 ;
        RECT 60.610 16.280 61.575 18.395 ;
        RECT 59.510 6.480 61.575 16.280 ;
        RECT 59.510 6.380 59.740 6.480 ;
        RECT 58.480 5.420 59.480 6.220 ;
        RECT 53.345 4.420 59.480 5.420 ;
      LAYER via ;
        RECT 136.060 205.300 137.060 206.300 ;
        RECT 139.760 205.430 140.760 206.430 ;
        RECT 151.540 202.370 152.540 203.370 ;
        RECT 81.080 200.610 81.380 200.910 ;
        RECT 143.440 201.200 144.440 202.200 ;
        RECT 105.820 200.530 106.120 200.830 ;
        RECT 129.070 200.520 129.370 200.820 ;
        RECT 152.700 200.510 153.000 200.810 ;
        RECT 59.600 198.310 60.800 199.510 ;
        RECT 71.400 198.960 72.400 199.220 ;
        RECT 59.490 194.800 60.460 195.800 ;
        RECT 6.855 188.260 7.865 189.270 ;
        RECT 59.540 186.735 60.550 187.745 ;
        RECT 64.100 184.770 64.400 186.630 ;
        RECT 70.790 198.490 71.050 198.760 ;
        RECT 65.700 198.030 70.110 198.300 ;
        RECT 65.660 197.390 69.430 197.660 ;
        RECT 66.340 196.750 70.110 197.020 ;
        RECT 65.660 196.110 69.430 196.380 ;
        RECT 66.340 195.470 70.110 195.740 ;
        RECT 65.660 194.830 69.430 195.100 ;
        RECT 66.340 194.190 70.110 194.460 ;
        RECT 65.660 193.550 69.430 193.820 ;
        RECT 66.340 192.910 70.110 193.180 ;
        RECT 65.660 192.270 69.430 192.540 ;
        RECT 66.340 191.630 70.110 191.900 ;
        RECT 65.660 190.990 69.430 191.260 ;
        RECT 66.340 190.350 70.110 190.620 ;
        RECT 65.660 189.710 69.430 189.980 ;
        RECT 66.340 189.070 70.110 189.340 ;
        RECT 65.660 188.430 69.430 188.700 ;
        RECT 66.340 187.790 70.110 188.060 ;
        RECT 65.660 187.150 69.430 187.420 ;
        RECT 66.340 186.510 70.110 186.780 ;
        RECT 65.660 185.870 69.430 186.140 ;
        RECT 66.340 185.230 70.110 185.500 ;
        RECT 71.400 198.030 72.400 198.290 ;
        RECT 73.630 198.960 75.080 199.220 ;
        RECT 73.630 198.490 75.080 198.760 ;
        RECT 73.630 198.030 75.080 198.290 ;
        RECT 76.150 198.900 76.450 199.190 ;
        RECT 77.480 198.440 78.920 198.700 ;
        RECT 77.480 198.030 78.920 198.290 ;
        RECT 80.200 198.410 81.200 199.410 ;
        RECT 71.400 196.860 72.400 197.120 ;
        RECT 71.400 195.930 72.400 196.190 ;
        RECT 73.630 196.860 75.080 197.120 ;
        RECT 73.630 196.390 75.080 196.660 ;
        RECT 73.630 195.930 75.080 196.190 ;
        RECT 76.170 197.330 76.430 197.600 ;
        RECT 77.480 196.860 78.920 197.120 ;
        RECT 77.480 196.450 78.920 196.710 ;
        RECT 80.200 196.860 81.200 197.120 ;
        RECT 65.660 184.590 70.110 184.860 ;
        RECT 76.170 193.490 76.430 193.760 ;
        RECT 74.080 193.010 78.520 193.280 ;
        RECT 74.080 192.370 78.520 192.640 ;
        RECT 74.080 191.730 78.520 192.000 ;
        RECT 74.080 191.090 78.520 191.360 ;
        RECT 74.080 190.450 78.520 190.720 ;
        RECT 74.080 189.810 78.520 190.080 ;
        RECT 74.080 189.170 78.520 189.440 ;
        RECT 74.080 188.530 78.520 188.800 ;
        RECT 71.400 182.410 72.400 183.410 ;
        RECT 84.340 198.230 85.540 199.430 ;
        RECT 96.140 198.880 97.140 199.140 ;
        RECT 84.280 186.655 85.290 187.665 ;
        RECT 88.840 184.690 89.140 186.550 ;
        RECT 95.530 198.410 95.790 198.680 ;
        RECT 90.440 197.950 94.850 198.220 ;
        RECT 90.400 197.310 94.170 197.580 ;
        RECT 91.080 196.670 94.850 196.940 ;
        RECT 90.400 196.030 94.170 196.300 ;
        RECT 91.080 195.390 94.850 195.660 ;
        RECT 90.400 194.750 94.170 195.020 ;
        RECT 91.080 194.110 94.850 194.380 ;
        RECT 90.400 193.470 94.170 193.740 ;
        RECT 91.080 192.830 94.850 193.100 ;
        RECT 90.400 192.190 94.170 192.460 ;
        RECT 91.080 191.550 94.850 191.820 ;
        RECT 90.400 190.910 94.170 191.180 ;
        RECT 91.080 190.270 94.850 190.540 ;
        RECT 90.400 189.630 94.170 189.900 ;
        RECT 91.080 188.990 94.850 189.260 ;
        RECT 90.400 188.350 94.170 188.620 ;
        RECT 91.080 187.710 94.850 187.980 ;
        RECT 90.400 187.070 94.170 187.340 ;
        RECT 91.080 186.430 94.850 186.700 ;
        RECT 90.400 185.790 94.170 186.060 ;
        RECT 91.080 185.150 94.850 185.420 ;
        RECT 96.140 197.950 97.140 198.210 ;
        RECT 98.370 198.880 99.820 199.140 ;
        RECT 98.370 198.410 99.820 198.680 ;
        RECT 98.370 197.950 99.820 198.210 ;
        RECT 100.890 198.820 101.190 199.110 ;
        RECT 102.220 198.360 103.660 198.620 ;
        RECT 102.220 197.950 103.660 198.210 ;
        RECT 104.940 198.330 105.940 199.330 ;
        RECT 96.140 196.780 97.140 197.040 ;
        RECT 96.140 195.850 97.140 196.110 ;
        RECT 98.370 196.780 99.820 197.040 ;
        RECT 98.370 196.310 99.820 196.580 ;
        RECT 98.370 195.850 99.820 196.110 ;
        RECT 100.910 197.250 101.170 197.520 ;
        RECT 102.220 196.780 103.660 197.040 ;
        RECT 102.220 196.370 103.660 196.630 ;
        RECT 104.940 196.780 105.940 197.040 ;
        RECT 90.400 184.510 94.850 184.780 ;
        RECT 100.910 193.410 101.170 193.680 ;
        RECT 98.820 192.930 103.260 193.200 ;
        RECT 98.820 192.290 103.260 192.560 ;
        RECT 98.820 191.650 103.260 191.920 ;
        RECT 98.820 191.010 103.260 191.280 ;
        RECT 98.820 190.370 103.260 190.640 ;
        RECT 98.820 189.730 103.260 190.000 ;
        RECT 98.820 189.090 103.260 189.360 ;
        RECT 98.820 188.450 103.260 188.720 ;
        RECT 96.140 182.330 97.140 183.330 ;
        RECT 107.590 198.220 108.790 199.420 ;
        RECT 119.390 198.870 120.390 199.130 ;
        RECT 107.530 186.645 108.540 187.655 ;
        RECT 112.090 184.680 112.390 186.540 ;
        RECT 118.780 198.400 119.040 198.670 ;
        RECT 113.690 197.940 118.100 198.210 ;
        RECT 113.650 197.300 117.420 197.570 ;
        RECT 114.330 196.660 118.100 196.930 ;
        RECT 113.650 196.020 117.420 196.290 ;
        RECT 114.330 195.380 118.100 195.650 ;
        RECT 113.650 194.740 117.420 195.010 ;
        RECT 114.330 194.100 118.100 194.370 ;
        RECT 113.650 193.460 117.420 193.730 ;
        RECT 114.330 192.820 118.100 193.090 ;
        RECT 113.650 192.180 117.420 192.450 ;
        RECT 114.330 191.540 118.100 191.810 ;
        RECT 113.650 190.900 117.420 191.170 ;
        RECT 114.330 190.260 118.100 190.530 ;
        RECT 113.650 189.620 117.420 189.890 ;
        RECT 114.330 188.980 118.100 189.250 ;
        RECT 113.650 188.340 117.420 188.610 ;
        RECT 114.330 187.700 118.100 187.970 ;
        RECT 113.650 187.060 117.420 187.330 ;
        RECT 114.330 186.420 118.100 186.690 ;
        RECT 113.650 185.780 117.420 186.050 ;
        RECT 114.330 185.140 118.100 185.410 ;
        RECT 119.390 197.940 120.390 198.200 ;
        RECT 121.620 198.870 123.070 199.130 ;
        RECT 121.620 198.400 123.070 198.670 ;
        RECT 121.620 197.940 123.070 198.200 ;
        RECT 124.140 198.810 124.440 199.100 ;
        RECT 125.470 198.350 126.910 198.610 ;
        RECT 125.470 197.940 126.910 198.200 ;
        RECT 128.190 198.320 129.190 199.320 ;
        RECT 119.390 196.770 120.390 197.030 ;
        RECT 119.390 195.840 120.390 196.100 ;
        RECT 121.620 196.770 123.070 197.030 ;
        RECT 121.620 196.300 123.070 196.570 ;
        RECT 121.620 195.840 123.070 196.100 ;
        RECT 124.160 197.240 124.420 197.510 ;
        RECT 125.470 196.770 126.910 197.030 ;
        RECT 125.470 196.360 126.910 196.620 ;
        RECT 128.190 196.770 129.190 197.030 ;
        RECT 113.650 184.500 118.100 184.770 ;
        RECT 124.160 193.400 124.420 193.670 ;
        RECT 122.070 192.920 126.510 193.190 ;
        RECT 122.070 192.280 126.510 192.550 ;
        RECT 122.070 191.640 126.510 191.910 ;
        RECT 122.070 191.000 126.510 191.270 ;
        RECT 122.070 190.360 126.510 190.630 ;
        RECT 122.070 189.720 126.510 189.990 ;
        RECT 122.070 189.080 126.510 189.350 ;
        RECT 122.070 188.440 126.510 188.710 ;
        RECT 119.390 182.320 120.390 183.320 ;
        RECT 131.220 198.210 132.420 199.410 ;
        RECT 143.020 198.860 144.020 199.120 ;
        RECT 131.160 186.635 132.170 187.645 ;
        RECT 135.720 184.670 136.020 186.530 ;
        RECT 142.410 198.390 142.670 198.660 ;
        RECT 137.320 197.930 141.730 198.200 ;
        RECT 137.280 197.290 141.050 197.560 ;
        RECT 137.960 196.650 141.730 196.920 ;
        RECT 137.280 196.010 141.050 196.280 ;
        RECT 137.960 195.370 141.730 195.640 ;
        RECT 137.280 194.730 141.050 195.000 ;
        RECT 137.960 194.090 141.730 194.360 ;
        RECT 137.280 193.450 141.050 193.720 ;
        RECT 137.960 192.810 141.730 193.080 ;
        RECT 137.280 192.170 141.050 192.440 ;
        RECT 137.960 191.530 141.730 191.800 ;
        RECT 137.280 190.890 141.050 191.160 ;
        RECT 137.960 190.250 141.730 190.520 ;
        RECT 137.280 189.610 141.050 189.880 ;
        RECT 137.960 188.970 141.730 189.240 ;
        RECT 137.280 188.330 141.050 188.600 ;
        RECT 137.960 187.690 141.730 187.960 ;
        RECT 137.280 187.050 141.050 187.320 ;
        RECT 137.960 186.410 141.730 186.680 ;
        RECT 137.280 185.770 141.050 186.040 ;
        RECT 137.960 185.130 141.730 185.400 ;
        RECT 143.020 197.930 144.020 198.190 ;
        RECT 145.250 198.860 146.700 199.120 ;
        RECT 145.250 198.390 146.700 198.660 ;
        RECT 145.250 197.930 146.700 198.190 ;
        RECT 147.770 198.800 148.070 199.090 ;
        RECT 149.100 198.340 150.540 198.600 ;
        RECT 149.100 197.930 150.540 198.190 ;
        RECT 151.820 198.310 152.820 199.310 ;
        RECT 143.020 196.760 144.020 197.020 ;
        RECT 143.020 195.830 144.020 196.090 ;
        RECT 145.250 196.760 146.700 197.020 ;
        RECT 145.250 196.290 146.700 196.560 ;
        RECT 145.250 195.830 146.700 196.090 ;
        RECT 147.790 197.230 148.050 197.500 ;
        RECT 149.100 196.760 150.540 197.020 ;
        RECT 149.100 196.350 150.540 196.610 ;
        RECT 151.820 196.760 152.820 197.020 ;
        RECT 137.280 184.490 141.730 184.760 ;
        RECT 147.790 193.390 148.050 193.660 ;
        RECT 145.700 192.910 150.140 193.180 ;
        RECT 145.700 192.270 150.140 192.540 ;
        RECT 145.700 191.630 150.140 191.900 ;
        RECT 145.700 190.990 150.140 191.260 ;
        RECT 145.700 190.350 150.140 190.620 ;
        RECT 145.700 189.710 150.140 189.980 ;
        RECT 145.700 189.070 150.140 189.340 ;
        RECT 145.700 188.430 150.140 188.700 ;
        RECT 143.020 182.310 144.020 183.310 ;
        RECT 72.750 180.590 73.750 181.590 ;
        RECT 97.490 180.510 98.490 181.510 ;
        RECT 120.740 180.500 121.740 181.500 ;
        RECT 144.370 180.490 145.370 181.490 ;
        RECT 151.860 180.520 152.860 181.520 ;
        RECT 80.970 174.520 81.270 174.820 ;
        RECT 104.150 174.430 104.450 174.730 ;
        RECT 127.050 174.630 127.350 174.930 ;
        RECT 150.150 174.740 150.450 175.040 ;
        RECT 59.490 172.220 60.690 173.420 ;
        RECT 71.290 172.870 72.290 173.130 ;
        RECT 46.990 167.030 47.990 168.030 ;
        RECT 8.205 162.445 9.215 163.455 ;
        RECT 59.430 160.645 60.440 161.655 ;
        RECT 63.990 158.680 64.290 160.540 ;
        RECT 70.680 172.400 70.940 172.670 ;
        RECT 65.590 171.940 70.000 172.210 ;
        RECT 65.550 171.300 69.320 171.570 ;
        RECT 66.230 170.660 70.000 170.930 ;
        RECT 65.550 170.020 69.320 170.290 ;
        RECT 66.230 169.380 70.000 169.650 ;
        RECT 65.550 168.740 69.320 169.010 ;
        RECT 66.230 168.100 70.000 168.370 ;
        RECT 65.550 167.460 69.320 167.730 ;
        RECT 66.230 166.820 70.000 167.090 ;
        RECT 65.550 166.180 69.320 166.450 ;
        RECT 66.230 165.540 70.000 165.810 ;
        RECT 65.550 164.900 69.320 165.170 ;
        RECT 66.230 164.260 70.000 164.530 ;
        RECT 65.550 163.620 69.320 163.890 ;
        RECT 66.230 162.980 70.000 163.250 ;
        RECT 65.550 162.340 69.320 162.610 ;
        RECT 66.230 161.700 70.000 161.970 ;
        RECT 65.550 161.060 69.320 161.330 ;
        RECT 66.230 160.420 70.000 160.690 ;
        RECT 65.550 159.780 69.320 160.050 ;
        RECT 66.230 159.140 70.000 159.410 ;
        RECT 71.290 171.940 72.290 172.200 ;
        RECT 73.520 172.870 74.970 173.130 ;
        RECT 73.520 172.400 74.970 172.670 ;
        RECT 73.520 171.940 74.970 172.200 ;
        RECT 76.040 172.810 76.340 173.100 ;
        RECT 77.370 172.350 78.810 172.610 ;
        RECT 77.370 171.940 78.810 172.200 ;
        RECT 80.090 172.320 81.090 173.320 ;
        RECT 71.290 170.770 72.290 171.030 ;
        RECT 71.290 169.840 72.290 170.100 ;
        RECT 73.520 170.770 74.970 171.030 ;
        RECT 73.520 170.300 74.970 170.570 ;
        RECT 73.520 169.840 74.970 170.100 ;
        RECT 76.060 171.240 76.320 171.510 ;
        RECT 77.370 170.770 78.810 171.030 ;
        RECT 77.370 170.360 78.810 170.620 ;
        RECT 80.090 170.770 81.090 171.030 ;
        RECT 65.550 158.500 70.000 158.770 ;
        RECT 76.060 167.400 76.320 167.670 ;
        RECT 73.970 166.920 78.410 167.190 ;
        RECT 73.970 166.280 78.410 166.550 ;
        RECT 73.970 165.640 78.410 165.910 ;
        RECT 73.970 165.000 78.410 165.270 ;
        RECT 73.970 164.360 78.410 164.630 ;
        RECT 73.970 163.720 78.410 163.990 ;
        RECT 73.970 163.080 78.410 163.350 ;
        RECT 73.970 162.440 78.410 162.710 ;
        RECT 71.290 156.320 72.290 157.320 ;
        RECT 82.670 172.130 83.870 173.330 ;
        RECT 94.470 172.780 95.470 173.040 ;
        RECT 82.610 160.555 83.620 161.565 ;
        RECT 87.170 158.590 87.470 160.450 ;
        RECT 93.860 172.310 94.120 172.580 ;
        RECT 88.770 171.850 93.180 172.120 ;
        RECT 88.730 171.210 92.500 171.480 ;
        RECT 89.410 170.570 93.180 170.840 ;
        RECT 88.730 169.930 92.500 170.200 ;
        RECT 89.410 169.290 93.180 169.560 ;
        RECT 88.730 168.650 92.500 168.920 ;
        RECT 89.410 168.010 93.180 168.280 ;
        RECT 88.730 167.370 92.500 167.640 ;
        RECT 89.410 166.730 93.180 167.000 ;
        RECT 88.730 166.090 92.500 166.360 ;
        RECT 89.410 165.450 93.180 165.720 ;
        RECT 88.730 164.810 92.500 165.080 ;
        RECT 89.410 164.170 93.180 164.440 ;
        RECT 88.730 163.530 92.500 163.800 ;
        RECT 89.410 162.890 93.180 163.160 ;
        RECT 88.730 162.250 92.500 162.520 ;
        RECT 89.410 161.610 93.180 161.880 ;
        RECT 88.730 160.970 92.500 161.240 ;
        RECT 89.410 160.330 93.180 160.600 ;
        RECT 88.730 159.690 92.500 159.960 ;
        RECT 89.410 159.050 93.180 159.320 ;
        RECT 94.470 171.850 95.470 172.110 ;
        RECT 96.700 172.780 98.150 173.040 ;
        RECT 96.700 172.310 98.150 172.580 ;
        RECT 96.700 171.850 98.150 172.110 ;
        RECT 99.220 172.720 99.520 173.010 ;
        RECT 100.550 172.260 101.990 172.520 ;
        RECT 100.550 171.850 101.990 172.110 ;
        RECT 103.270 172.230 104.270 173.230 ;
        RECT 94.470 170.680 95.470 170.940 ;
        RECT 94.470 169.750 95.470 170.010 ;
        RECT 96.700 170.680 98.150 170.940 ;
        RECT 96.700 170.210 98.150 170.480 ;
        RECT 96.700 169.750 98.150 170.010 ;
        RECT 99.240 171.150 99.500 171.420 ;
        RECT 100.550 170.680 101.990 170.940 ;
        RECT 100.550 170.270 101.990 170.530 ;
        RECT 103.270 170.680 104.270 170.940 ;
        RECT 88.730 158.410 93.180 158.680 ;
        RECT 99.240 167.310 99.500 167.580 ;
        RECT 97.150 166.830 101.590 167.100 ;
        RECT 97.150 166.190 101.590 166.460 ;
        RECT 97.150 165.550 101.590 165.820 ;
        RECT 97.150 164.910 101.590 165.180 ;
        RECT 97.150 164.270 101.590 164.540 ;
        RECT 97.150 163.630 101.590 163.900 ;
        RECT 97.150 162.990 101.590 163.260 ;
        RECT 97.150 162.350 101.590 162.620 ;
        RECT 94.470 156.230 95.470 157.230 ;
        RECT 105.570 172.330 106.770 173.530 ;
        RECT 117.370 172.980 118.370 173.240 ;
        RECT 105.510 160.755 106.520 161.765 ;
        RECT 110.070 158.790 110.370 160.650 ;
        RECT 116.760 172.510 117.020 172.780 ;
        RECT 111.670 172.050 116.080 172.320 ;
        RECT 111.630 171.410 115.400 171.680 ;
        RECT 112.310 170.770 116.080 171.040 ;
        RECT 111.630 170.130 115.400 170.400 ;
        RECT 112.310 169.490 116.080 169.760 ;
        RECT 111.630 168.850 115.400 169.120 ;
        RECT 112.310 168.210 116.080 168.480 ;
        RECT 111.630 167.570 115.400 167.840 ;
        RECT 112.310 166.930 116.080 167.200 ;
        RECT 111.630 166.290 115.400 166.560 ;
        RECT 112.310 165.650 116.080 165.920 ;
        RECT 111.630 165.010 115.400 165.280 ;
        RECT 112.310 164.370 116.080 164.640 ;
        RECT 111.630 163.730 115.400 164.000 ;
        RECT 112.310 163.090 116.080 163.360 ;
        RECT 111.630 162.450 115.400 162.720 ;
        RECT 112.310 161.810 116.080 162.080 ;
        RECT 111.630 161.170 115.400 161.440 ;
        RECT 112.310 160.530 116.080 160.800 ;
        RECT 111.630 159.890 115.400 160.160 ;
        RECT 112.310 159.250 116.080 159.520 ;
        RECT 117.370 172.050 118.370 172.310 ;
        RECT 119.600 172.980 121.050 173.240 ;
        RECT 119.600 172.510 121.050 172.780 ;
        RECT 119.600 172.050 121.050 172.310 ;
        RECT 122.120 172.920 122.420 173.210 ;
        RECT 123.450 172.460 124.890 172.720 ;
        RECT 123.450 172.050 124.890 172.310 ;
        RECT 126.170 172.430 127.170 173.430 ;
        RECT 117.370 170.880 118.370 171.140 ;
        RECT 117.370 169.950 118.370 170.210 ;
        RECT 119.600 170.880 121.050 171.140 ;
        RECT 119.600 170.410 121.050 170.680 ;
        RECT 119.600 169.950 121.050 170.210 ;
        RECT 122.140 171.350 122.400 171.620 ;
        RECT 123.450 170.880 124.890 171.140 ;
        RECT 123.450 170.470 124.890 170.730 ;
        RECT 126.170 170.880 127.170 171.140 ;
        RECT 111.630 158.610 116.080 158.880 ;
        RECT 122.140 167.510 122.400 167.780 ;
        RECT 120.050 167.030 124.490 167.300 ;
        RECT 120.050 166.390 124.490 166.660 ;
        RECT 120.050 165.750 124.490 166.020 ;
        RECT 120.050 165.110 124.490 165.380 ;
        RECT 120.050 164.470 124.490 164.740 ;
        RECT 120.050 163.830 124.490 164.100 ;
        RECT 120.050 163.190 124.490 163.460 ;
        RECT 120.050 162.550 124.490 162.820 ;
        RECT 117.370 156.430 118.370 157.430 ;
        RECT 128.670 172.440 129.870 173.640 ;
        RECT 140.470 173.090 141.470 173.350 ;
        RECT 128.610 160.865 129.620 161.875 ;
        RECT 133.170 158.900 133.470 160.760 ;
        RECT 139.860 172.620 140.120 172.890 ;
        RECT 134.770 172.160 139.180 172.430 ;
        RECT 134.730 171.520 138.500 171.790 ;
        RECT 135.410 170.880 139.180 171.150 ;
        RECT 134.730 170.240 138.500 170.510 ;
        RECT 135.410 169.600 139.180 169.870 ;
        RECT 134.730 168.960 138.500 169.230 ;
        RECT 135.410 168.320 139.180 168.590 ;
        RECT 134.730 167.680 138.500 167.950 ;
        RECT 135.410 167.040 139.180 167.310 ;
        RECT 134.730 166.400 138.500 166.670 ;
        RECT 135.410 165.760 139.180 166.030 ;
        RECT 134.730 165.120 138.500 165.390 ;
        RECT 135.410 164.480 139.180 164.750 ;
        RECT 134.730 163.840 138.500 164.110 ;
        RECT 135.410 163.200 139.180 163.470 ;
        RECT 134.730 162.560 138.500 162.830 ;
        RECT 135.410 161.920 139.180 162.190 ;
        RECT 134.730 161.280 138.500 161.550 ;
        RECT 135.410 160.640 139.180 160.910 ;
        RECT 134.730 160.000 138.500 160.270 ;
        RECT 135.410 159.360 139.180 159.630 ;
        RECT 140.470 172.160 141.470 172.420 ;
        RECT 142.700 173.090 144.150 173.350 ;
        RECT 142.700 172.620 144.150 172.890 ;
        RECT 142.700 172.160 144.150 172.420 ;
        RECT 145.220 173.030 145.520 173.320 ;
        RECT 146.550 172.570 147.990 172.830 ;
        RECT 146.550 172.160 147.990 172.420 ;
        RECT 149.270 172.540 150.270 173.540 ;
        RECT 140.470 170.990 141.470 171.250 ;
        RECT 140.470 170.060 141.470 170.320 ;
        RECT 142.700 170.990 144.150 171.250 ;
        RECT 142.700 170.520 144.150 170.790 ;
        RECT 142.700 170.060 144.150 170.320 ;
        RECT 145.240 171.460 145.500 171.730 ;
        RECT 146.550 170.990 147.990 171.250 ;
        RECT 146.550 170.580 147.990 170.840 ;
        RECT 149.270 170.990 150.270 171.250 ;
        RECT 134.730 158.720 139.180 158.990 ;
        RECT 145.240 167.620 145.500 167.890 ;
        RECT 143.150 167.140 147.590 167.410 ;
        RECT 143.150 166.500 147.590 166.770 ;
        RECT 143.150 165.860 147.590 166.130 ;
        RECT 143.150 165.220 147.590 165.490 ;
        RECT 143.150 164.580 147.590 164.850 ;
        RECT 143.150 163.940 147.590 164.210 ;
        RECT 143.150 163.300 147.590 163.570 ;
        RECT 143.150 162.660 147.590 162.930 ;
        RECT 140.470 156.540 141.470 157.540 ;
        RECT 72.640 154.500 73.640 155.500 ;
        RECT 95.820 154.410 96.820 155.410 ;
        RECT 118.720 154.610 119.720 155.610 ;
        RECT 141.820 154.720 142.820 155.720 ;
        RECT 104.360 148.790 104.660 149.090 ;
        RECT 127.390 148.940 127.690 149.240 ;
        RECT 150.400 149.020 150.700 149.320 ;
        RECT 82.880 146.490 84.080 147.690 ;
        RECT 94.680 147.140 95.680 147.400 ;
        RECT 57.170 141.310 58.170 142.310 ;
        RECT 8.265 136.770 9.275 137.780 ;
        RECT 82.820 134.915 83.830 135.925 ;
        RECT 87.380 132.950 87.680 134.810 ;
        RECT 94.070 146.670 94.330 146.940 ;
        RECT 88.980 146.210 93.390 146.480 ;
        RECT 88.940 145.570 92.710 145.840 ;
        RECT 89.620 144.930 93.390 145.200 ;
        RECT 88.940 144.290 92.710 144.560 ;
        RECT 89.620 143.650 93.390 143.920 ;
        RECT 88.940 143.010 92.710 143.280 ;
        RECT 89.620 142.370 93.390 142.640 ;
        RECT 88.940 141.730 92.710 142.000 ;
        RECT 89.620 141.090 93.390 141.360 ;
        RECT 88.940 140.450 92.710 140.720 ;
        RECT 89.620 139.810 93.390 140.080 ;
        RECT 88.940 139.170 92.710 139.440 ;
        RECT 89.620 138.530 93.390 138.800 ;
        RECT 88.940 137.890 92.710 138.160 ;
        RECT 89.620 137.250 93.390 137.520 ;
        RECT 88.940 136.610 92.710 136.880 ;
        RECT 89.620 135.970 93.390 136.240 ;
        RECT 88.940 135.330 92.710 135.600 ;
        RECT 89.620 134.690 93.390 134.960 ;
        RECT 88.940 134.050 92.710 134.320 ;
        RECT 89.620 133.410 93.390 133.680 ;
        RECT 94.680 146.210 95.680 146.470 ;
        RECT 96.910 147.140 98.360 147.400 ;
        RECT 96.910 146.670 98.360 146.940 ;
        RECT 96.910 146.210 98.360 146.470 ;
        RECT 99.430 147.080 99.730 147.370 ;
        RECT 100.760 146.620 102.200 146.880 ;
        RECT 100.760 146.210 102.200 146.470 ;
        RECT 103.480 146.590 104.480 147.590 ;
        RECT 94.680 145.040 95.680 145.300 ;
        RECT 94.680 144.110 95.680 144.370 ;
        RECT 96.910 145.040 98.360 145.300 ;
        RECT 96.910 144.570 98.360 144.840 ;
        RECT 96.910 144.110 98.360 144.370 ;
        RECT 99.450 145.510 99.710 145.780 ;
        RECT 100.760 145.040 102.200 145.300 ;
        RECT 100.760 144.630 102.200 144.890 ;
        RECT 103.480 145.040 104.480 145.300 ;
        RECT 88.940 132.770 93.390 133.040 ;
        RECT 99.450 141.670 99.710 141.940 ;
        RECT 97.360 141.190 101.800 141.460 ;
        RECT 97.360 140.550 101.800 140.820 ;
        RECT 97.360 139.910 101.800 140.180 ;
        RECT 97.360 139.270 101.800 139.540 ;
        RECT 97.360 138.630 101.800 138.900 ;
        RECT 97.360 137.990 101.800 138.260 ;
        RECT 97.360 137.350 101.800 137.620 ;
        RECT 97.360 136.710 101.800 136.980 ;
        RECT 94.680 130.590 95.680 131.590 ;
        RECT 105.910 146.640 107.110 147.840 ;
        RECT 117.710 147.290 118.710 147.550 ;
        RECT 105.850 135.065 106.860 136.075 ;
        RECT 110.410 133.100 110.710 134.960 ;
        RECT 117.100 146.820 117.360 147.090 ;
        RECT 112.010 146.360 116.420 146.630 ;
        RECT 111.970 145.720 115.740 145.990 ;
        RECT 112.650 145.080 116.420 145.350 ;
        RECT 111.970 144.440 115.740 144.710 ;
        RECT 112.650 143.800 116.420 144.070 ;
        RECT 111.970 143.160 115.740 143.430 ;
        RECT 112.650 142.520 116.420 142.790 ;
        RECT 111.970 141.880 115.740 142.150 ;
        RECT 112.650 141.240 116.420 141.510 ;
        RECT 111.970 140.600 115.740 140.870 ;
        RECT 112.650 139.960 116.420 140.230 ;
        RECT 111.970 139.320 115.740 139.590 ;
        RECT 112.650 138.680 116.420 138.950 ;
        RECT 111.970 138.040 115.740 138.310 ;
        RECT 112.650 137.400 116.420 137.670 ;
        RECT 111.970 136.760 115.740 137.030 ;
        RECT 112.650 136.120 116.420 136.390 ;
        RECT 111.970 135.480 115.740 135.750 ;
        RECT 112.650 134.840 116.420 135.110 ;
        RECT 111.970 134.200 115.740 134.470 ;
        RECT 112.650 133.560 116.420 133.830 ;
        RECT 117.710 146.360 118.710 146.620 ;
        RECT 119.940 147.290 121.390 147.550 ;
        RECT 119.940 146.820 121.390 147.090 ;
        RECT 119.940 146.360 121.390 146.620 ;
        RECT 122.460 147.230 122.760 147.520 ;
        RECT 123.790 146.770 125.230 147.030 ;
        RECT 123.790 146.360 125.230 146.620 ;
        RECT 126.510 146.740 127.510 147.740 ;
        RECT 117.710 145.190 118.710 145.450 ;
        RECT 117.710 144.260 118.710 144.520 ;
        RECT 119.940 145.190 121.390 145.450 ;
        RECT 119.940 144.720 121.390 144.990 ;
        RECT 119.940 144.260 121.390 144.520 ;
        RECT 122.480 145.660 122.740 145.930 ;
        RECT 123.790 145.190 125.230 145.450 ;
        RECT 123.790 144.780 125.230 145.040 ;
        RECT 126.510 145.190 127.510 145.450 ;
        RECT 111.970 132.920 116.420 133.190 ;
        RECT 122.480 141.820 122.740 142.090 ;
        RECT 120.390 141.340 124.830 141.610 ;
        RECT 120.390 140.700 124.830 140.970 ;
        RECT 120.390 140.060 124.830 140.330 ;
        RECT 120.390 139.420 124.830 139.690 ;
        RECT 120.390 138.780 124.830 139.050 ;
        RECT 120.390 138.140 124.830 138.410 ;
        RECT 120.390 137.500 124.830 137.770 ;
        RECT 120.390 136.860 124.830 137.130 ;
        RECT 117.710 130.740 118.710 131.740 ;
        RECT 128.920 146.720 130.120 147.920 ;
        RECT 140.720 147.370 141.720 147.630 ;
        RECT 128.860 135.145 129.870 136.155 ;
        RECT 133.420 133.180 133.720 135.040 ;
        RECT 140.110 146.900 140.370 147.170 ;
        RECT 135.020 146.440 139.430 146.710 ;
        RECT 134.980 145.800 138.750 146.070 ;
        RECT 135.660 145.160 139.430 145.430 ;
        RECT 134.980 144.520 138.750 144.790 ;
        RECT 135.660 143.880 139.430 144.150 ;
        RECT 134.980 143.240 138.750 143.510 ;
        RECT 135.660 142.600 139.430 142.870 ;
        RECT 134.980 141.960 138.750 142.230 ;
        RECT 135.660 141.320 139.430 141.590 ;
        RECT 134.980 140.680 138.750 140.950 ;
        RECT 135.660 140.040 139.430 140.310 ;
        RECT 134.980 139.400 138.750 139.670 ;
        RECT 135.660 138.760 139.430 139.030 ;
        RECT 134.980 138.120 138.750 138.390 ;
        RECT 135.660 137.480 139.430 137.750 ;
        RECT 134.980 136.840 138.750 137.110 ;
        RECT 135.660 136.200 139.430 136.470 ;
        RECT 134.980 135.560 138.750 135.830 ;
        RECT 135.660 134.920 139.430 135.190 ;
        RECT 134.980 134.280 138.750 134.550 ;
        RECT 135.660 133.640 139.430 133.910 ;
        RECT 140.720 146.440 141.720 146.700 ;
        RECT 142.950 147.370 144.400 147.630 ;
        RECT 142.950 146.900 144.400 147.170 ;
        RECT 142.950 146.440 144.400 146.700 ;
        RECT 145.470 147.310 145.770 147.600 ;
        RECT 146.800 146.850 148.240 147.110 ;
        RECT 146.800 146.440 148.240 146.700 ;
        RECT 149.520 146.820 150.520 147.820 ;
        RECT 140.720 145.270 141.720 145.530 ;
        RECT 140.720 144.340 141.720 144.600 ;
        RECT 142.950 145.270 144.400 145.530 ;
        RECT 142.950 144.800 144.400 145.070 ;
        RECT 142.950 144.340 144.400 144.600 ;
        RECT 145.490 145.740 145.750 146.010 ;
        RECT 146.800 145.270 148.240 145.530 ;
        RECT 146.800 144.860 148.240 145.120 ;
        RECT 149.520 145.270 150.520 145.530 ;
        RECT 134.980 133.000 139.430 133.270 ;
        RECT 145.490 141.900 145.750 142.170 ;
        RECT 143.400 141.420 147.840 141.690 ;
        RECT 143.400 140.780 147.840 141.050 ;
        RECT 143.400 140.140 147.840 140.410 ;
        RECT 143.400 139.500 147.840 139.770 ;
        RECT 143.400 138.860 147.840 139.130 ;
        RECT 143.400 138.220 147.840 138.490 ;
        RECT 143.400 137.580 147.840 137.850 ;
        RECT 143.400 136.940 147.840 137.210 ;
        RECT 140.720 130.820 141.720 131.820 ;
        RECT 96.030 128.770 97.030 129.770 ;
        RECT 119.060 128.920 120.060 129.920 ;
        RECT 142.070 129.000 143.070 130.000 ;
        RECT 55.480 28.140 56.980 29.640 ;
        RECT 51.275 19.165 52.600 20.490 ;
        RECT 60.395 19.135 61.765 20.505 ;
        RECT 55.610 10.560 57.110 12.060 ;
      LAYER met2 ;
        RECT 136.060 206.300 137.060 207.785 ;
        RECT 139.760 206.430 140.760 208.125 ;
        RECT 136.030 205.300 137.090 206.300 ;
        RECT 139.730 205.430 140.790 206.430 ;
        RECT 143.440 201.170 144.440 205.105 ;
        RECT 151.540 203.370 152.540 205.305 ;
        RECT 151.510 202.370 152.570 203.370 ;
        RECT 81.850 200.910 82.130 200.945 ;
        RECT 81.050 200.610 82.140 200.910 ;
        RECT 106.590 200.830 106.870 200.865 ;
        RECT 81.850 200.575 82.130 200.610 ;
        RECT 105.790 200.530 106.880 200.830 ;
        RECT 129.840 200.820 130.120 200.855 ;
        RECT 106.590 200.495 106.870 200.530 ;
        RECT 129.040 200.520 130.130 200.820 ;
        RECT 153.470 200.810 153.750 200.845 ;
        RECT 129.840 200.485 130.120 200.520 ;
        RECT 152.670 200.510 153.760 200.810 ;
        RECT 153.470 200.475 153.750 200.510 ;
        RECT 59.600 199.485 60.800 199.540 ;
        RECT 59.580 198.335 60.820 199.485 ;
        RECT 71.300 198.960 75.110 199.220 ;
        RECT 76.100 198.900 76.500 199.190 ;
        RECT 70.760 198.490 76.400 198.760 ;
        RECT 80.100 198.700 81.300 199.510 ;
        RECT 84.340 199.405 85.540 199.460 ;
        RECT 59.600 198.280 60.800 198.335 ;
        RECT 65.630 198.030 70.140 198.300 ;
        RECT 76.200 198.290 76.400 198.490 ;
        RECT 77.450 198.440 81.300 198.700 ;
        RECT 80.100 198.310 81.300 198.440 ;
        RECT 71.300 198.030 75.110 198.290 ;
        RECT 76.200 198.030 78.950 198.290 ;
        RECT 84.320 198.255 85.560 199.405 ;
        RECT 96.040 198.880 99.850 199.140 ;
        RECT 100.840 198.820 101.240 199.110 ;
        RECT 95.500 198.410 101.140 198.680 ;
        RECT 104.840 198.620 106.040 199.430 ;
        RECT 107.590 199.395 108.790 199.450 ;
        RECT 84.340 198.200 85.540 198.255 ;
        RECT 64.970 197.390 69.460 197.660 ;
        RECT 64.970 196.380 65.970 197.390 ;
        RECT 69.800 197.020 70.800 198.030 ;
        RECT 76.200 197.630 76.400 198.030 ;
        RECT 90.370 197.950 94.880 198.220 ;
        RECT 100.940 198.210 101.140 198.410 ;
        RECT 102.190 198.360 106.040 198.620 ;
        RECT 104.840 198.230 106.040 198.360 ;
        RECT 107.570 198.245 108.810 199.395 ;
        RECT 119.290 198.870 123.100 199.130 ;
        RECT 124.090 198.810 124.490 199.100 ;
        RECT 118.750 198.400 124.390 198.670 ;
        RECT 128.090 198.610 129.290 199.420 ;
        RECT 131.220 199.385 132.420 199.440 ;
        RECT 96.040 197.950 99.850 198.210 ;
        RECT 100.940 197.950 103.690 198.210 ;
        RECT 107.590 198.190 108.790 198.245 ;
        RECT 76.170 197.300 76.430 197.630 ;
        RECT 89.710 197.310 94.200 197.580 ;
        RECT 66.310 196.750 70.800 197.020 ;
        RECT 71.300 196.860 75.110 197.120 ;
        RECT 77.450 196.860 81.300 197.120 ;
        RECT 64.970 196.110 69.460 196.380 ;
        RECT 46.620 193.800 47.620 195.255 ;
        RECT 59.490 194.770 60.460 195.830 ;
        RECT 64.970 195.100 65.970 196.110 ;
        RECT 69.800 195.740 70.800 196.750 ;
        RECT 76.200 196.660 78.950 196.710 ;
        RECT 73.600 196.450 78.950 196.660 ;
        RECT 73.600 196.390 76.400 196.450 ;
        RECT 71.300 195.930 75.110 196.190 ;
        RECT 66.310 195.470 70.800 195.740 ;
        RECT 64.970 194.830 69.460 195.100 ;
        RECT 64.970 193.820 65.970 194.830 ;
        RECT 69.800 194.460 70.800 195.470 ;
        RECT 66.310 194.190 70.800 194.460 ;
        RECT 46.590 192.800 47.650 193.800 ;
        RECT 64.970 193.550 69.460 193.820 ;
        RECT 64.970 192.820 65.970 193.550 ;
        RECT 69.800 193.180 70.800 194.190 ;
        RECT 76.200 193.790 76.400 196.390 ;
        RECT 89.710 196.300 90.710 197.310 ;
        RECT 94.540 196.940 95.540 197.950 ;
        RECT 100.940 197.550 101.140 197.950 ;
        RECT 113.620 197.940 118.130 198.210 ;
        RECT 124.190 198.200 124.390 198.400 ;
        RECT 125.440 198.350 129.290 198.610 ;
        RECT 128.090 198.220 129.290 198.350 ;
        RECT 131.200 198.235 132.440 199.385 ;
        RECT 142.920 198.860 146.730 199.120 ;
        RECT 147.720 198.800 148.120 199.090 ;
        RECT 142.380 198.390 148.020 198.660 ;
        RECT 151.720 198.600 152.920 199.410 ;
        RECT 119.290 197.940 123.100 198.200 ;
        RECT 124.190 197.940 126.940 198.200 ;
        RECT 131.220 198.180 132.420 198.235 ;
        RECT 100.910 197.220 101.170 197.550 ;
        RECT 112.960 197.300 117.450 197.570 ;
        RECT 91.050 196.670 95.540 196.940 ;
        RECT 96.040 196.780 99.850 197.040 ;
        RECT 102.190 196.780 106.040 197.040 ;
        RECT 89.710 196.030 94.200 196.300 ;
        RECT 89.710 195.020 90.710 196.030 ;
        RECT 94.540 195.660 95.540 196.670 ;
        RECT 100.940 196.580 103.690 196.630 ;
        RECT 98.340 196.370 103.690 196.580 ;
        RECT 98.340 196.310 101.140 196.370 ;
        RECT 96.040 195.850 99.850 196.110 ;
        RECT 91.050 195.390 95.540 195.660 ;
        RECT 89.710 194.750 94.200 195.020 ;
        RECT 76.170 193.460 76.430 193.790 ;
        RECT 89.710 193.740 90.710 194.750 ;
        RECT 94.540 194.380 95.540 195.390 ;
        RECT 91.050 194.110 95.540 194.380 ;
        RECT 89.710 193.470 94.200 193.740 ;
        RECT 66.310 192.910 70.800 193.180 ;
        RECT 74.050 193.010 79.850 193.280 ;
        RECT 63.970 192.540 65.970 192.820 ;
        RECT 63.970 192.270 69.460 192.540 ;
        RECT 63.970 191.260 65.970 192.270 ;
        RECT 69.800 191.910 70.800 192.910 ;
        RECT 72.750 192.370 78.550 192.640 ;
        RECT 72.750 191.910 73.750 192.370 ;
        RECT 78.850 192.000 79.850 193.010 ;
        RECT 89.710 192.740 90.710 193.470 ;
        RECT 94.540 193.100 95.540 194.110 ;
        RECT 100.940 193.710 101.140 196.310 ;
        RECT 112.960 196.290 113.960 197.300 ;
        RECT 117.790 196.930 118.790 197.940 ;
        RECT 124.190 197.540 124.390 197.940 ;
        RECT 137.250 197.930 141.760 198.200 ;
        RECT 147.820 198.190 148.020 198.390 ;
        RECT 149.070 198.340 152.920 198.600 ;
        RECT 151.720 198.210 152.920 198.340 ;
        RECT 142.920 197.930 146.730 198.190 ;
        RECT 147.820 197.930 150.570 198.190 ;
        RECT 124.160 197.210 124.420 197.540 ;
        RECT 136.590 197.290 141.080 197.560 ;
        RECT 114.300 196.660 118.790 196.930 ;
        RECT 119.290 196.770 123.100 197.030 ;
        RECT 125.440 196.770 129.290 197.030 ;
        RECT 112.960 196.020 117.450 196.290 ;
        RECT 112.960 195.010 113.960 196.020 ;
        RECT 117.790 195.650 118.790 196.660 ;
        RECT 124.190 196.570 126.940 196.620 ;
        RECT 121.590 196.360 126.940 196.570 ;
        RECT 121.590 196.300 124.390 196.360 ;
        RECT 119.290 195.840 123.100 196.100 ;
        RECT 114.300 195.380 118.790 195.650 ;
        RECT 112.960 194.740 117.450 195.010 ;
        RECT 112.960 193.730 113.960 194.740 ;
        RECT 117.790 194.370 118.790 195.380 ;
        RECT 114.300 194.100 118.790 194.370 ;
        RECT 100.910 193.380 101.170 193.710 ;
        RECT 112.960 193.460 117.450 193.730 ;
        RECT 91.050 192.830 95.540 193.100 ;
        RECT 98.790 192.930 104.590 193.200 ;
        RECT 69.800 191.900 73.750 191.910 ;
        RECT 66.310 191.630 73.750 191.900 ;
        RECT 74.050 191.860 79.850 192.000 ;
        RECT 88.710 192.460 90.710 192.740 ;
        RECT 88.710 192.190 94.200 192.460 ;
        RECT 74.050 191.730 81.300 191.860 ;
        RECT 69.800 191.360 73.750 191.630 ;
        RECT 63.970 190.990 69.460 191.260 ;
        RECT 69.800 191.090 78.550 191.360 ;
        RECT 63.970 189.980 65.970 190.990 ;
        RECT 69.800 190.620 73.750 191.090 ;
        RECT 78.850 190.720 81.300 191.730 ;
        RECT 66.310 190.350 73.750 190.620 ;
        RECT 74.050 190.450 81.300 190.720 ;
        RECT 69.800 190.080 73.750 190.350 ;
        RECT 63.970 189.710 69.460 189.980 ;
        RECT 69.800 189.910 78.550 190.080 ;
        RECT 4.235 189.270 5.245 189.315 ;
        RECT 6.855 189.270 7.865 189.300 ;
        RECT 4.235 188.260 7.865 189.270 ;
        RECT 4.235 188.215 5.245 188.260 ;
        RECT 6.855 188.230 7.865 188.260 ;
        RECT 63.970 188.700 65.970 189.710 ;
        RECT 69.800 189.340 70.800 189.910 ;
        RECT 66.310 189.070 70.800 189.340 ;
        RECT 63.970 188.430 69.460 188.700 ;
        RECT 59.510 186.735 60.580 187.745 ;
        RECT 63.970 187.420 65.970 188.430 ;
        RECT 69.800 188.060 70.800 189.070 ;
        RECT 66.310 187.790 70.800 188.060 ;
        RECT 63.970 187.150 69.460 187.420 ;
        RECT 59.540 185.460 60.550 186.735 ;
        RECT 63.970 186.140 65.970 187.150 ;
        RECT 69.800 186.780 70.800 187.790 ;
        RECT 66.310 186.510 70.800 186.780 ;
        RECT 63.970 185.870 69.460 186.140 ;
        RECT 63.970 184.860 65.970 185.870 ;
        RECT 69.800 185.500 70.800 186.510 ;
        RECT 72.750 189.810 78.550 189.910 ;
        RECT 78.850 189.860 81.300 190.450 ;
        RECT 88.710 191.180 90.710 192.190 ;
        RECT 94.540 191.830 95.540 192.830 ;
        RECT 97.490 192.290 103.290 192.560 ;
        RECT 97.490 191.830 98.490 192.290 ;
        RECT 103.590 191.920 104.590 192.930 ;
        RECT 112.960 192.730 113.960 193.460 ;
        RECT 117.790 193.090 118.790 194.100 ;
        RECT 124.190 193.700 124.390 196.300 ;
        RECT 136.590 196.280 137.590 197.290 ;
        RECT 141.420 196.920 142.420 197.930 ;
        RECT 147.820 197.530 148.020 197.930 ;
        RECT 147.790 197.200 148.050 197.530 ;
        RECT 137.930 196.650 142.420 196.920 ;
        RECT 142.920 196.760 146.730 197.020 ;
        RECT 149.070 196.760 152.920 197.020 ;
        RECT 136.590 196.010 141.080 196.280 ;
        RECT 136.590 195.000 137.590 196.010 ;
        RECT 141.420 195.640 142.420 196.650 ;
        RECT 147.820 196.560 150.570 196.610 ;
        RECT 145.220 196.350 150.570 196.560 ;
        RECT 145.220 196.290 148.020 196.350 ;
        RECT 142.920 195.830 146.730 196.090 ;
        RECT 137.930 195.370 142.420 195.640 ;
        RECT 136.590 194.730 141.080 195.000 ;
        RECT 136.590 193.720 137.590 194.730 ;
        RECT 141.420 194.360 142.420 195.370 ;
        RECT 137.930 194.090 142.420 194.360 ;
        RECT 124.160 193.370 124.420 193.700 ;
        RECT 136.590 193.450 141.080 193.720 ;
        RECT 114.300 192.820 118.790 193.090 ;
        RECT 122.040 192.920 127.840 193.190 ;
        RECT 94.540 191.820 98.490 191.830 ;
        RECT 91.050 191.550 98.490 191.820 ;
        RECT 98.790 191.780 104.590 191.920 ;
        RECT 111.960 192.450 113.960 192.730 ;
        RECT 111.960 192.180 117.450 192.450 ;
        RECT 98.790 191.650 106.040 191.780 ;
        RECT 94.540 191.280 98.490 191.550 ;
        RECT 88.710 190.910 94.200 191.180 ;
        RECT 94.540 191.010 103.290 191.280 ;
        RECT 88.710 189.900 90.710 190.910 ;
        RECT 94.540 190.540 98.490 191.010 ;
        RECT 103.590 190.640 106.040 191.650 ;
        RECT 91.050 190.270 98.490 190.540 ;
        RECT 98.790 190.370 106.040 190.640 ;
        RECT 94.540 190.000 98.490 190.270 ;
        RECT 72.750 188.800 73.750 189.810 ;
        RECT 78.850 189.440 79.850 189.860 ;
        RECT 74.050 189.170 79.850 189.440 ;
        RECT 79.670 189.160 79.850 189.170 ;
        RECT 88.710 189.630 94.200 189.900 ;
        RECT 94.540 189.830 103.290 190.000 ;
        RECT 72.750 188.530 78.550 188.800 ;
        RECT 88.710 188.620 90.710 189.630 ;
        RECT 94.540 189.260 95.540 189.830 ;
        RECT 91.050 188.990 95.540 189.260 ;
        RECT 66.310 185.230 70.140 185.500 ;
        RECT 69.800 185.220 70.140 185.230 ;
        RECT 63.970 182.860 70.420 184.860 ;
        RECT 71.300 182.310 72.500 183.510 ;
        RECT 72.750 180.560 73.750 188.530 ;
        RECT 88.710 188.350 94.200 188.620 ;
        RECT 84.250 186.655 85.320 187.665 ;
        RECT 88.710 187.340 90.710 188.350 ;
        RECT 94.540 187.980 95.540 188.990 ;
        RECT 91.050 187.710 95.540 187.980 ;
        RECT 88.710 187.070 94.200 187.340 ;
        RECT 84.280 185.380 85.290 186.655 ;
        RECT 88.710 186.060 90.710 187.070 ;
        RECT 94.540 186.700 95.540 187.710 ;
        RECT 91.050 186.430 95.540 186.700 ;
        RECT 88.710 185.790 94.200 186.060 ;
        RECT 88.710 184.780 90.710 185.790 ;
        RECT 94.540 185.420 95.540 186.430 ;
        RECT 97.490 189.730 103.290 189.830 ;
        RECT 103.590 189.780 106.040 190.370 ;
        RECT 111.960 191.170 113.960 192.180 ;
        RECT 117.790 191.820 118.790 192.820 ;
        RECT 120.740 192.280 126.540 192.550 ;
        RECT 120.740 191.820 121.740 192.280 ;
        RECT 126.840 191.910 127.840 192.920 ;
        RECT 136.590 192.720 137.590 193.450 ;
        RECT 141.420 193.080 142.420 194.090 ;
        RECT 147.820 193.690 148.020 196.290 ;
        RECT 147.790 193.360 148.050 193.690 ;
        RECT 137.930 192.810 142.420 193.080 ;
        RECT 145.670 192.910 151.470 193.180 ;
        RECT 117.790 191.810 121.740 191.820 ;
        RECT 114.300 191.540 121.740 191.810 ;
        RECT 122.040 191.770 127.840 191.910 ;
        RECT 135.590 192.440 137.590 192.720 ;
        RECT 135.590 192.170 141.080 192.440 ;
        RECT 122.040 191.640 129.290 191.770 ;
        RECT 117.790 191.270 121.740 191.540 ;
        RECT 111.960 190.900 117.450 191.170 ;
        RECT 117.790 191.000 126.540 191.270 ;
        RECT 111.960 189.890 113.960 190.900 ;
        RECT 117.790 190.530 121.740 191.000 ;
        RECT 126.840 190.630 129.290 191.640 ;
        RECT 114.300 190.260 121.740 190.530 ;
        RECT 122.040 190.360 129.290 190.630 ;
        RECT 117.790 189.990 121.740 190.260 ;
        RECT 97.490 188.720 98.490 189.730 ;
        RECT 103.590 189.360 104.590 189.780 ;
        RECT 98.790 189.090 104.590 189.360 ;
        RECT 104.410 189.080 104.590 189.090 ;
        RECT 111.960 189.620 117.450 189.890 ;
        RECT 117.790 189.820 126.540 189.990 ;
        RECT 97.490 188.450 103.290 188.720 ;
        RECT 111.960 188.610 113.960 189.620 ;
        RECT 117.790 189.250 118.790 189.820 ;
        RECT 114.300 188.980 118.790 189.250 ;
        RECT 91.050 185.150 94.880 185.420 ;
        RECT 94.540 185.140 94.880 185.150 ;
        RECT 88.710 182.780 95.160 184.780 ;
        RECT 96.040 182.230 97.240 183.430 ;
        RECT 97.490 180.480 98.490 188.450 ;
        RECT 111.960 188.340 117.450 188.610 ;
        RECT 107.500 186.645 108.570 187.655 ;
        RECT 111.960 187.330 113.960 188.340 ;
        RECT 117.790 187.970 118.790 188.980 ;
        RECT 114.300 187.700 118.790 187.970 ;
        RECT 111.960 187.060 117.450 187.330 ;
        RECT 107.530 185.370 108.540 186.645 ;
        RECT 111.960 186.050 113.960 187.060 ;
        RECT 117.790 186.690 118.790 187.700 ;
        RECT 114.300 186.420 118.790 186.690 ;
        RECT 111.960 185.780 117.450 186.050 ;
        RECT 111.960 184.770 113.960 185.780 ;
        RECT 117.790 185.410 118.790 186.420 ;
        RECT 120.740 189.720 126.540 189.820 ;
        RECT 126.840 189.770 129.290 190.360 ;
        RECT 135.590 191.160 137.590 192.170 ;
        RECT 141.420 191.810 142.420 192.810 ;
        RECT 144.370 192.270 150.170 192.540 ;
        RECT 144.370 191.810 145.370 192.270 ;
        RECT 150.470 191.900 151.470 192.910 ;
        RECT 141.420 191.800 145.370 191.810 ;
        RECT 137.930 191.530 145.370 191.800 ;
        RECT 145.670 191.760 151.470 191.900 ;
        RECT 145.670 191.630 152.920 191.760 ;
        RECT 141.420 191.260 145.370 191.530 ;
        RECT 135.590 190.890 141.080 191.160 ;
        RECT 141.420 190.990 150.170 191.260 ;
        RECT 135.590 189.880 137.590 190.890 ;
        RECT 141.420 190.520 145.370 190.990 ;
        RECT 150.470 190.620 152.920 191.630 ;
        RECT 137.930 190.250 145.370 190.520 ;
        RECT 145.670 190.350 152.920 190.620 ;
        RECT 141.420 189.980 145.370 190.250 ;
        RECT 120.740 188.710 121.740 189.720 ;
        RECT 126.840 189.350 127.840 189.770 ;
        RECT 122.040 189.080 127.840 189.350 ;
        RECT 127.660 189.070 127.840 189.080 ;
        RECT 135.590 189.610 141.080 189.880 ;
        RECT 141.420 189.810 150.170 189.980 ;
        RECT 120.740 188.440 126.540 188.710 ;
        RECT 135.590 188.600 137.590 189.610 ;
        RECT 141.420 189.240 142.420 189.810 ;
        RECT 137.930 188.970 142.420 189.240 ;
        RECT 114.300 185.140 118.130 185.410 ;
        RECT 117.790 185.130 118.130 185.140 ;
        RECT 111.960 182.770 118.410 184.770 ;
        RECT 119.290 182.220 120.490 183.420 ;
        RECT 120.740 180.470 121.740 188.440 ;
        RECT 135.590 188.330 141.080 188.600 ;
        RECT 131.130 186.635 132.200 187.645 ;
        RECT 135.590 187.320 137.590 188.330 ;
        RECT 141.420 187.960 142.420 188.970 ;
        RECT 137.930 187.690 142.420 187.960 ;
        RECT 135.590 187.050 141.080 187.320 ;
        RECT 131.160 185.360 132.170 186.635 ;
        RECT 135.590 186.040 137.590 187.050 ;
        RECT 141.420 186.680 142.420 187.690 ;
        RECT 137.930 186.410 142.420 186.680 ;
        RECT 135.590 185.770 141.080 186.040 ;
        RECT 135.590 184.760 137.590 185.770 ;
        RECT 141.420 185.400 142.420 186.410 ;
        RECT 144.370 189.710 150.170 189.810 ;
        RECT 150.470 189.760 152.920 190.350 ;
        RECT 144.370 188.700 145.370 189.710 ;
        RECT 150.470 189.340 151.470 189.760 ;
        RECT 145.670 189.070 151.470 189.340 ;
        RECT 151.290 189.060 151.470 189.070 ;
        RECT 144.370 188.430 150.170 188.700 ;
        RECT 137.930 185.130 141.760 185.400 ;
        RECT 141.420 185.120 141.760 185.130 ;
        RECT 135.590 182.760 142.040 184.760 ;
        RECT 142.920 182.210 144.120 183.410 ;
        RECT 144.370 180.460 145.370 188.430 ;
        RECT 151.860 179.385 152.860 181.550 ;
        RECT 150.920 175.040 151.200 175.075 ;
        RECT 127.820 174.930 128.100 174.965 ;
        RECT 81.740 174.820 82.020 174.855 ;
        RECT 80.940 174.520 82.030 174.820 ;
        RECT 104.920 174.730 105.200 174.765 ;
        RECT 81.740 174.485 82.020 174.520 ;
        RECT 104.120 174.430 105.210 174.730 ;
        RECT 127.020 174.630 128.110 174.930 ;
        RECT 150.120 174.740 151.210 175.040 ;
        RECT 150.920 174.705 151.200 174.740 ;
        RECT 127.820 174.595 128.100 174.630 ;
        RECT 104.920 174.395 105.200 174.430 ;
        RECT 127.775 173.960 128.145 174.240 ;
        RECT 128.670 173.615 129.870 173.670 ;
        RECT 105.570 173.505 106.770 173.560 ;
        RECT 59.490 173.395 60.690 173.450 ;
        RECT 59.470 172.245 60.710 173.395 ;
        RECT 71.190 172.870 75.000 173.130 ;
        RECT 75.990 172.810 76.390 173.100 ;
        RECT 70.650 172.400 76.290 172.670 ;
        RECT 79.990 172.610 81.190 173.420 ;
        RECT 82.670 173.305 83.870 173.360 ;
        RECT 59.490 172.190 60.690 172.245 ;
        RECT 65.520 171.940 70.030 172.210 ;
        RECT 76.090 172.200 76.290 172.400 ;
        RECT 77.340 172.350 81.190 172.610 ;
        RECT 79.990 172.220 81.190 172.350 ;
        RECT 71.190 171.940 75.000 172.200 ;
        RECT 76.090 171.940 78.840 172.200 ;
        RECT 82.650 172.155 83.890 173.305 ;
        RECT 94.370 172.780 98.180 173.040 ;
        RECT 99.170 172.720 99.570 173.010 ;
        RECT 93.830 172.310 99.470 172.580 ;
        RECT 103.170 172.520 104.370 173.330 ;
        RECT 82.670 172.100 83.870 172.155 ;
        RECT 64.860 171.300 69.350 171.570 ;
        RECT 64.860 170.290 65.860 171.300 ;
        RECT 69.690 170.930 70.690 171.940 ;
        RECT 76.090 171.540 76.290 171.940 ;
        RECT 88.700 171.850 93.210 172.120 ;
        RECT 99.270 172.110 99.470 172.310 ;
        RECT 100.520 172.260 104.370 172.520 ;
        RECT 105.550 172.355 106.790 173.505 ;
        RECT 117.270 172.980 121.080 173.240 ;
        RECT 122.070 172.920 122.470 173.210 ;
        RECT 116.730 172.510 122.370 172.780 ;
        RECT 126.070 172.720 127.270 173.530 ;
        RECT 105.570 172.300 106.770 172.355 ;
        RECT 103.170 172.130 104.370 172.260 ;
        RECT 94.370 171.850 98.180 172.110 ;
        RECT 99.270 171.850 102.020 172.110 ;
        RECT 111.600 172.050 116.110 172.320 ;
        RECT 122.170 172.310 122.370 172.510 ;
        RECT 123.420 172.460 127.270 172.720 ;
        RECT 128.650 172.465 129.890 173.615 ;
        RECT 140.370 173.090 144.180 173.350 ;
        RECT 145.170 173.030 145.570 173.320 ;
        RECT 139.830 172.620 145.470 172.890 ;
        RECT 149.170 172.830 150.370 173.640 ;
        RECT 126.070 172.330 127.270 172.460 ;
        RECT 128.670 172.410 129.870 172.465 ;
        RECT 117.270 172.050 121.080 172.310 ;
        RECT 122.170 172.050 124.920 172.310 ;
        RECT 134.700 172.160 139.210 172.430 ;
        RECT 145.270 172.420 145.470 172.620 ;
        RECT 146.520 172.570 150.370 172.830 ;
        RECT 149.170 172.440 150.370 172.570 ;
        RECT 140.370 172.160 144.180 172.420 ;
        RECT 145.270 172.160 148.020 172.420 ;
        RECT 76.060 171.210 76.320 171.540 ;
        RECT 88.040 171.210 92.530 171.480 ;
        RECT 66.200 170.660 70.690 170.930 ;
        RECT 71.190 170.770 75.000 171.030 ;
        RECT 77.340 170.770 81.190 171.030 ;
        RECT 64.860 170.020 69.350 170.290 ;
        RECT 46.990 167.000 47.990 169.435 ;
        RECT 64.860 169.010 65.860 170.020 ;
        RECT 69.690 169.650 70.690 170.660 ;
        RECT 76.090 170.570 78.840 170.620 ;
        RECT 73.490 170.360 78.840 170.570 ;
        RECT 73.490 170.300 76.290 170.360 ;
        RECT 71.190 169.840 75.000 170.100 ;
        RECT 66.200 169.380 70.690 169.650 ;
        RECT 64.860 168.740 69.350 169.010 ;
        RECT 64.860 167.730 65.860 168.740 ;
        RECT 69.690 168.370 70.690 169.380 ;
        RECT 66.200 168.100 70.690 168.370 ;
        RECT 64.860 167.460 69.350 167.730 ;
        RECT 64.860 166.730 65.860 167.460 ;
        RECT 69.690 167.090 70.690 168.100 ;
        RECT 76.090 167.700 76.290 170.300 ;
        RECT 88.040 170.200 89.040 171.210 ;
        RECT 92.870 170.840 93.870 171.850 ;
        RECT 99.270 171.450 99.470 171.850 ;
        RECT 99.240 171.120 99.500 171.450 ;
        RECT 110.940 171.410 115.430 171.680 ;
        RECT 89.380 170.570 93.870 170.840 ;
        RECT 94.370 170.680 98.180 170.940 ;
        RECT 100.520 170.680 104.370 170.940 ;
        RECT 88.040 169.930 92.530 170.200 ;
        RECT 88.040 168.920 89.040 169.930 ;
        RECT 92.870 169.560 93.870 170.570 ;
        RECT 99.270 170.480 102.020 170.530 ;
        RECT 96.670 170.270 102.020 170.480 ;
        RECT 110.940 170.400 111.940 171.410 ;
        RECT 115.770 171.040 116.770 172.050 ;
        RECT 122.170 171.650 122.370 172.050 ;
        RECT 122.140 171.320 122.400 171.650 ;
        RECT 134.040 171.520 138.530 171.790 ;
        RECT 112.280 170.770 116.770 171.040 ;
        RECT 117.270 170.880 121.080 171.140 ;
        RECT 123.420 170.880 127.270 171.140 ;
        RECT 96.670 170.210 99.470 170.270 ;
        RECT 94.370 169.750 98.180 170.010 ;
        RECT 89.380 169.290 93.870 169.560 ;
        RECT 88.040 168.650 92.530 168.920 ;
        RECT 76.060 167.370 76.320 167.700 ;
        RECT 88.040 167.640 89.040 168.650 ;
        RECT 92.870 168.280 93.870 169.290 ;
        RECT 89.380 168.010 93.870 168.280 ;
        RECT 88.040 167.370 92.530 167.640 ;
        RECT 66.200 166.820 70.690 167.090 ;
        RECT 73.940 166.920 79.740 167.190 ;
        RECT 63.860 166.450 65.860 166.730 ;
        RECT 63.860 166.180 69.350 166.450 ;
        RECT 63.860 165.170 65.860 166.180 ;
        RECT 69.690 165.820 70.690 166.820 ;
        RECT 72.640 166.280 78.440 166.550 ;
        RECT 72.640 165.820 73.640 166.280 ;
        RECT 78.740 165.910 79.740 166.920 ;
        RECT 88.040 166.640 89.040 167.370 ;
        RECT 92.870 167.000 93.870 168.010 ;
        RECT 99.270 167.610 99.470 170.210 ;
        RECT 110.940 170.130 115.430 170.400 ;
        RECT 110.940 169.120 111.940 170.130 ;
        RECT 115.770 169.760 116.770 170.770 ;
        RECT 122.170 170.680 124.920 170.730 ;
        RECT 119.570 170.470 124.920 170.680 ;
        RECT 134.040 170.510 135.040 171.520 ;
        RECT 138.870 171.150 139.870 172.160 ;
        RECT 145.270 171.760 145.470 172.160 ;
        RECT 145.240 171.430 145.500 171.760 ;
        RECT 135.380 170.880 139.870 171.150 ;
        RECT 140.370 170.990 144.180 171.250 ;
        RECT 146.520 170.990 150.370 171.250 ;
        RECT 119.570 170.410 122.370 170.470 ;
        RECT 117.270 169.950 121.080 170.210 ;
        RECT 112.280 169.490 116.770 169.760 ;
        RECT 110.940 168.850 115.430 169.120 ;
        RECT 110.940 167.840 111.940 168.850 ;
        RECT 115.770 168.480 116.770 169.490 ;
        RECT 112.280 168.210 116.770 168.480 ;
        RECT 99.240 167.280 99.500 167.610 ;
        RECT 110.940 167.570 115.430 167.840 ;
        RECT 89.380 166.730 93.870 167.000 ;
        RECT 97.120 166.830 102.920 167.100 ;
        RECT 110.940 166.840 111.940 167.570 ;
        RECT 115.770 167.200 116.770 168.210 ;
        RECT 122.170 167.810 122.370 170.410 ;
        RECT 134.040 170.240 138.530 170.510 ;
        RECT 134.040 169.230 135.040 170.240 ;
        RECT 138.870 169.870 139.870 170.880 ;
        RECT 145.270 170.790 148.020 170.840 ;
        RECT 142.670 170.580 148.020 170.790 ;
        RECT 142.670 170.520 145.470 170.580 ;
        RECT 140.370 170.060 144.180 170.320 ;
        RECT 135.380 169.600 139.870 169.870 ;
        RECT 134.040 168.960 138.530 169.230 ;
        RECT 134.040 167.950 135.040 168.960 ;
        RECT 138.870 168.590 139.870 169.600 ;
        RECT 135.380 168.320 139.870 168.590 ;
        RECT 122.140 167.480 122.400 167.810 ;
        RECT 134.040 167.680 138.530 167.950 ;
        RECT 112.280 166.930 116.770 167.200 ;
        RECT 120.020 167.030 125.820 167.300 ;
        RECT 69.690 165.810 73.640 165.820 ;
        RECT 66.200 165.540 73.640 165.810 ;
        RECT 73.940 165.770 79.740 165.910 ;
        RECT 87.040 166.360 89.040 166.640 ;
        RECT 87.040 166.090 92.530 166.360 ;
        RECT 73.940 165.640 81.190 165.770 ;
        RECT 69.690 165.270 73.640 165.540 ;
        RECT 63.860 164.900 69.350 165.170 ;
        RECT 69.690 165.000 78.440 165.270 ;
        RECT 63.860 163.890 65.860 164.900 ;
        RECT 69.690 164.530 73.640 165.000 ;
        RECT 78.740 164.630 81.190 165.640 ;
        RECT 66.200 164.260 73.640 164.530 ;
        RECT 73.940 164.360 81.190 164.630 ;
        RECT 69.690 163.990 73.640 164.260 ;
        RECT 63.860 163.620 69.350 163.890 ;
        RECT 69.690 163.820 78.440 163.990 ;
        RECT 8.205 163.455 9.215 163.485 ;
        RECT 6.700 162.445 9.215 163.455 ;
        RECT 8.205 162.415 9.215 162.445 ;
        RECT 63.860 162.610 65.860 163.620 ;
        RECT 69.690 163.250 70.690 163.820 ;
        RECT 66.200 162.980 70.690 163.250 ;
        RECT 63.860 162.340 69.350 162.610 ;
        RECT 59.400 160.645 60.470 161.655 ;
        RECT 63.860 161.330 65.860 162.340 ;
        RECT 69.690 161.970 70.690 162.980 ;
        RECT 66.200 161.700 70.690 161.970 ;
        RECT 63.860 161.060 69.350 161.330 ;
        RECT 59.430 159.370 60.440 160.645 ;
        RECT 63.860 160.050 65.860 161.060 ;
        RECT 69.690 160.690 70.690 161.700 ;
        RECT 66.200 160.420 70.690 160.690 ;
        RECT 63.860 159.780 69.350 160.050 ;
        RECT 63.860 158.770 65.860 159.780 ;
        RECT 69.690 159.410 70.690 160.420 ;
        RECT 72.640 163.720 78.440 163.820 ;
        RECT 78.740 163.770 81.190 164.360 ;
        RECT 87.040 165.080 89.040 166.090 ;
        RECT 92.870 165.730 93.870 166.730 ;
        RECT 95.820 166.190 101.620 166.460 ;
        RECT 95.820 165.730 96.820 166.190 ;
        RECT 101.920 165.820 102.920 166.830 ;
        RECT 92.870 165.720 96.820 165.730 ;
        RECT 89.380 165.450 96.820 165.720 ;
        RECT 97.120 165.680 102.920 165.820 ;
        RECT 109.940 166.560 111.940 166.840 ;
        RECT 109.940 166.290 115.430 166.560 ;
        RECT 97.120 165.550 104.370 165.680 ;
        RECT 92.870 165.180 96.820 165.450 ;
        RECT 87.040 164.810 92.530 165.080 ;
        RECT 92.870 164.910 101.620 165.180 ;
        RECT 87.040 163.800 89.040 164.810 ;
        RECT 92.870 164.440 96.820 164.910 ;
        RECT 101.920 164.540 104.370 165.550 ;
        RECT 89.380 164.170 96.820 164.440 ;
        RECT 97.120 164.270 104.370 164.540 ;
        RECT 92.870 163.900 96.820 164.170 ;
        RECT 72.640 162.710 73.640 163.720 ;
        RECT 78.740 163.350 79.740 163.770 ;
        RECT 73.940 163.080 79.740 163.350 ;
        RECT 79.560 163.070 79.740 163.080 ;
        RECT 87.040 163.530 92.530 163.800 ;
        RECT 92.870 163.730 101.620 163.900 ;
        RECT 72.640 162.440 78.440 162.710 ;
        RECT 87.040 162.520 89.040 163.530 ;
        RECT 92.870 163.160 93.870 163.730 ;
        RECT 89.380 162.890 93.870 163.160 ;
        RECT 66.200 159.140 70.030 159.410 ;
        RECT 69.690 159.130 70.030 159.140 ;
        RECT 63.860 156.770 70.310 158.770 ;
        RECT 71.190 156.220 72.390 157.420 ;
        RECT 72.640 154.470 73.640 162.440 ;
        RECT 87.040 162.250 92.530 162.520 ;
        RECT 82.580 160.555 83.650 161.565 ;
        RECT 87.040 161.240 89.040 162.250 ;
        RECT 92.870 161.880 93.870 162.890 ;
        RECT 89.380 161.610 93.870 161.880 ;
        RECT 87.040 160.970 92.530 161.240 ;
        RECT 82.610 159.280 83.620 160.555 ;
        RECT 87.040 159.960 89.040 160.970 ;
        RECT 92.870 160.600 93.870 161.610 ;
        RECT 89.380 160.330 93.870 160.600 ;
        RECT 87.040 159.690 92.530 159.960 ;
        RECT 87.040 158.680 89.040 159.690 ;
        RECT 92.870 159.320 93.870 160.330 ;
        RECT 95.820 163.630 101.620 163.730 ;
        RECT 101.920 163.680 104.370 164.270 ;
        RECT 109.940 165.280 111.940 166.290 ;
        RECT 115.770 165.930 116.770 166.930 ;
        RECT 118.720 166.390 124.520 166.660 ;
        RECT 118.720 165.930 119.720 166.390 ;
        RECT 124.820 166.020 125.820 167.030 ;
        RECT 134.040 166.950 135.040 167.680 ;
        RECT 138.870 167.310 139.870 168.320 ;
        RECT 145.270 167.920 145.470 170.520 ;
        RECT 145.240 167.590 145.500 167.920 ;
        RECT 135.380 167.040 139.870 167.310 ;
        RECT 143.120 167.140 148.920 167.410 ;
        RECT 115.770 165.920 119.720 165.930 ;
        RECT 112.280 165.650 119.720 165.920 ;
        RECT 120.020 165.880 125.820 166.020 ;
        RECT 133.040 166.670 135.040 166.950 ;
        RECT 133.040 166.400 138.530 166.670 ;
        RECT 120.020 165.750 127.270 165.880 ;
        RECT 115.770 165.380 119.720 165.650 ;
        RECT 109.940 165.010 115.430 165.280 ;
        RECT 115.770 165.110 124.520 165.380 ;
        RECT 109.940 164.000 111.940 165.010 ;
        RECT 115.770 164.640 119.720 165.110 ;
        RECT 124.820 164.740 127.270 165.750 ;
        RECT 112.280 164.370 119.720 164.640 ;
        RECT 120.020 164.470 127.270 164.740 ;
        RECT 115.770 164.100 119.720 164.370 ;
        RECT 109.940 163.730 115.430 164.000 ;
        RECT 115.770 163.930 124.520 164.100 ;
        RECT 95.820 162.620 96.820 163.630 ;
        RECT 101.920 163.260 102.920 163.680 ;
        RECT 97.120 162.990 102.920 163.260 ;
        RECT 102.740 162.980 102.920 162.990 ;
        RECT 109.940 162.720 111.940 163.730 ;
        RECT 115.770 163.360 116.770 163.930 ;
        RECT 112.280 163.090 116.770 163.360 ;
        RECT 95.820 162.350 101.620 162.620 ;
        RECT 109.940 162.450 115.430 162.720 ;
        RECT 89.380 159.050 93.210 159.320 ;
        RECT 92.870 159.040 93.210 159.050 ;
        RECT 87.040 156.680 93.490 158.680 ;
        RECT 94.370 156.130 95.570 157.330 ;
        RECT 95.820 154.380 96.820 162.350 ;
        RECT 105.480 160.755 106.550 161.765 ;
        RECT 109.940 161.440 111.940 162.450 ;
        RECT 115.770 162.080 116.770 163.090 ;
        RECT 112.280 161.810 116.770 162.080 ;
        RECT 109.940 161.170 115.430 161.440 ;
        RECT 105.510 159.480 106.520 160.755 ;
        RECT 109.940 160.160 111.940 161.170 ;
        RECT 115.770 160.800 116.770 161.810 ;
        RECT 112.280 160.530 116.770 160.800 ;
        RECT 109.940 159.890 115.430 160.160 ;
        RECT 109.940 158.880 111.940 159.890 ;
        RECT 115.770 159.520 116.770 160.530 ;
        RECT 118.720 163.830 124.520 163.930 ;
        RECT 124.820 163.880 127.270 164.470 ;
        RECT 133.040 165.390 135.040 166.400 ;
        RECT 138.870 166.040 139.870 167.040 ;
        RECT 141.820 166.500 147.620 166.770 ;
        RECT 141.820 166.040 142.820 166.500 ;
        RECT 147.920 166.130 148.920 167.140 ;
        RECT 138.870 166.030 142.820 166.040 ;
        RECT 135.380 165.760 142.820 166.030 ;
        RECT 143.120 165.990 148.920 166.130 ;
        RECT 143.120 165.860 150.370 165.990 ;
        RECT 138.870 165.490 142.820 165.760 ;
        RECT 133.040 165.120 138.530 165.390 ;
        RECT 138.870 165.220 147.620 165.490 ;
        RECT 133.040 164.110 135.040 165.120 ;
        RECT 138.870 164.750 142.820 165.220 ;
        RECT 147.920 164.850 150.370 165.860 ;
        RECT 135.380 164.480 142.820 164.750 ;
        RECT 143.120 164.580 150.370 164.850 ;
        RECT 138.870 164.210 142.820 164.480 ;
        RECT 118.720 162.820 119.720 163.830 ;
        RECT 124.820 163.460 125.820 163.880 ;
        RECT 120.020 163.190 125.820 163.460 ;
        RECT 125.640 163.180 125.820 163.190 ;
        RECT 133.040 163.840 138.530 164.110 ;
        RECT 138.870 164.040 147.620 164.210 ;
        RECT 133.040 162.830 135.040 163.840 ;
        RECT 138.870 163.470 139.870 164.040 ;
        RECT 135.380 163.200 139.870 163.470 ;
        RECT 118.720 162.550 124.520 162.820 ;
        RECT 133.040 162.560 138.530 162.830 ;
        RECT 112.280 159.250 116.110 159.520 ;
        RECT 115.770 159.240 116.110 159.250 ;
        RECT 109.940 156.880 116.390 158.880 ;
        RECT 117.270 156.330 118.470 157.530 ;
        RECT 118.720 154.580 119.720 162.550 ;
        RECT 128.580 160.865 129.650 161.875 ;
        RECT 133.040 161.550 135.040 162.560 ;
        RECT 138.870 162.190 139.870 163.200 ;
        RECT 135.380 161.920 139.870 162.190 ;
        RECT 133.040 161.280 138.530 161.550 ;
        RECT 128.610 159.590 129.620 160.865 ;
        RECT 133.040 160.270 135.040 161.280 ;
        RECT 138.870 160.910 139.870 161.920 ;
        RECT 135.380 160.640 139.870 160.910 ;
        RECT 133.040 160.000 138.530 160.270 ;
        RECT 133.040 158.990 135.040 160.000 ;
        RECT 138.870 159.630 139.870 160.640 ;
        RECT 141.820 163.940 147.620 164.040 ;
        RECT 147.920 163.990 150.370 164.580 ;
        RECT 141.820 162.930 142.820 163.940 ;
        RECT 147.920 163.570 148.920 163.990 ;
        RECT 143.120 163.300 148.920 163.570 ;
        RECT 148.740 163.290 148.920 163.300 ;
        RECT 141.820 162.660 147.620 162.930 ;
        RECT 135.380 159.360 139.210 159.630 ;
        RECT 138.870 159.350 139.210 159.360 ;
        RECT 133.040 156.990 139.490 158.990 ;
        RECT 140.370 156.440 141.570 157.640 ;
        RECT 141.820 155.660 142.820 162.660 ;
        RECT 141.775 154.660 142.865 155.660 ;
        RECT 151.170 149.320 151.450 149.355 ;
        RECT 128.160 149.240 128.440 149.275 ;
        RECT 105.130 149.090 105.410 149.125 ;
        RECT 104.330 148.790 105.420 149.090 ;
        RECT 127.360 148.940 128.450 149.240 ;
        RECT 150.370 149.020 151.460 149.320 ;
        RECT 151.170 148.985 151.450 149.020 ;
        RECT 128.160 148.905 128.440 148.940 ;
        RECT 105.130 148.755 105.410 148.790 ;
        RECT 128.920 147.895 130.120 147.950 ;
        RECT 105.910 147.815 107.110 147.870 ;
        RECT 82.880 147.665 84.080 147.720 ;
        RECT 82.860 146.515 84.100 147.665 ;
        RECT 94.580 147.140 98.390 147.400 ;
        RECT 99.380 147.080 99.780 147.370 ;
        RECT 94.040 146.670 99.680 146.940 ;
        RECT 103.380 146.880 104.580 147.690 ;
        RECT 82.880 146.460 84.080 146.515 ;
        RECT 88.910 146.210 93.420 146.480 ;
        RECT 99.480 146.470 99.680 146.670 ;
        RECT 100.730 146.620 104.580 146.880 ;
        RECT 105.890 146.665 107.130 147.815 ;
        RECT 117.610 147.290 121.420 147.550 ;
        RECT 122.410 147.230 122.810 147.520 ;
        RECT 117.070 146.820 122.710 147.090 ;
        RECT 126.410 147.030 127.610 147.840 ;
        RECT 103.380 146.490 104.580 146.620 ;
        RECT 105.910 146.610 107.110 146.665 ;
        RECT 94.580 146.210 98.390 146.470 ;
        RECT 99.480 146.210 102.230 146.470 ;
        RECT 111.940 146.360 116.450 146.630 ;
        RECT 122.510 146.620 122.710 146.820 ;
        RECT 123.760 146.770 127.610 147.030 ;
        RECT 126.410 146.640 127.610 146.770 ;
        RECT 128.900 146.745 130.140 147.895 ;
        RECT 140.620 147.370 144.430 147.630 ;
        RECT 145.420 147.310 145.820 147.600 ;
        RECT 140.080 146.900 145.720 147.170 ;
        RECT 149.420 147.110 150.620 147.920 ;
        RECT 128.920 146.690 130.120 146.745 ;
        RECT 117.610 146.360 121.420 146.620 ;
        RECT 122.510 146.360 125.260 146.620 ;
        RECT 134.950 146.440 139.460 146.710 ;
        RECT 145.520 146.700 145.720 146.900 ;
        RECT 146.770 146.850 150.620 147.110 ;
        RECT 149.420 146.720 150.620 146.850 ;
        RECT 140.620 146.440 144.430 146.700 ;
        RECT 145.520 146.440 148.270 146.700 ;
        RECT 88.250 145.570 92.740 145.840 ;
        RECT 88.250 144.560 89.250 145.570 ;
        RECT 93.080 145.200 94.080 146.210 ;
        RECT 99.480 145.810 99.680 146.210 ;
        RECT 99.450 145.480 99.710 145.810 ;
        RECT 111.280 145.720 115.770 145.990 ;
        RECT 89.590 144.930 94.080 145.200 ;
        RECT 94.580 145.040 98.390 145.300 ;
        RECT 100.730 145.040 104.580 145.300 ;
        RECT 88.250 144.290 92.740 144.560 ;
        RECT 88.250 143.280 89.250 144.290 ;
        RECT 93.080 143.920 94.080 144.930 ;
        RECT 99.480 144.840 102.230 144.890 ;
        RECT 96.880 144.630 102.230 144.840 ;
        RECT 111.280 144.710 112.280 145.720 ;
        RECT 116.110 145.350 117.110 146.360 ;
        RECT 122.510 145.960 122.710 146.360 ;
        RECT 122.480 145.630 122.740 145.960 ;
        RECT 134.290 145.800 138.780 146.070 ;
        RECT 112.620 145.080 117.110 145.350 ;
        RECT 117.610 145.190 121.420 145.450 ;
        RECT 123.760 145.190 127.610 145.450 ;
        RECT 96.880 144.570 99.680 144.630 ;
        RECT 94.580 144.110 98.390 144.370 ;
        RECT 89.590 143.650 94.080 143.920 ;
        RECT 88.250 143.010 92.740 143.280 ;
        RECT 57.170 142.310 58.170 142.340 ;
        RECT 57.125 141.310 58.215 142.310 ;
        RECT 88.250 142.000 89.250 143.010 ;
        RECT 93.080 142.640 94.080 143.650 ;
        RECT 89.590 142.370 94.080 142.640 ;
        RECT 88.250 141.730 92.740 142.000 ;
        RECT 57.170 141.280 58.170 141.310 ;
        RECT 88.250 141.000 89.250 141.730 ;
        RECT 93.080 141.360 94.080 142.370 ;
        RECT 99.480 141.970 99.680 144.570 ;
        RECT 111.280 144.440 115.770 144.710 ;
        RECT 111.280 143.430 112.280 144.440 ;
        RECT 116.110 144.070 117.110 145.080 ;
        RECT 122.510 144.990 125.260 145.040 ;
        RECT 119.910 144.780 125.260 144.990 ;
        RECT 134.290 144.790 135.290 145.800 ;
        RECT 139.120 145.430 140.120 146.440 ;
        RECT 145.520 146.040 145.720 146.440 ;
        RECT 145.490 145.710 145.750 146.040 ;
        RECT 135.630 145.160 140.120 145.430 ;
        RECT 140.620 145.270 144.430 145.530 ;
        RECT 146.770 145.270 150.620 145.530 ;
        RECT 119.910 144.720 122.710 144.780 ;
        RECT 117.610 144.260 121.420 144.520 ;
        RECT 112.620 143.800 117.110 144.070 ;
        RECT 111.280 143.160 115.770 143.430 ;
        RECT 111.280 142.150 112.280 143.160 ;
        RECT 116.110 142.790 117.110 143.800 ;
        RECT 112.620 142.520 117.110 142.790 ;
        RECT 99.450 141.640 99.710 141.970 ;
        RECT 111.280 141.880 115.770 142.150 ;
        RECT 89.590 141.090 94.080 141.360 ;
        RECT 97.330 141.190 103.130 141.460 ;
        RECT 87.250 140.720 89.250 141.000 ;
        RECT 87.250 140.450 92.740 140.720 ;
        RECT 87.250 139.440 89.250 140.450 ;
        RECT 93.080 140.090 94.080 141.090 ;
        RECT 96.030 140.550 101.830 140.820 ;
        RECT 96.030 140.090 97.030 140.550 ;
        RECT 102.130 140.180 103.130 141.190 ;
        RECT 111.280 141.150 112.280 141.880 ;
        RECT 116.110 141.510 117.110 142.520 ;
        RECT 122.510 142.120 122.710 144.720 ;
        RECT 134.290 144.520 138.780 144.790 ;
        RECT 134.290 143.510 135.290 144.520 ;
        RECT 139.120 144.150 140.120 145.160 ;
        RECT 145.520 145.070 148.270 145.120 ;
        RECT 142.920 144.860 148.270 145.070 ;
        RECT 142.920 144.800 145.720 144.860 ;
        RECT 140.620 144.340 144.430 144.600 ;
        RECT 135.630 143.880 140.120 144.150 ;
        RECT 134.290 143.240 138.780 143.510 ;
        RECT 134.290 142.230 135.290 143.240 ;
        RECT 139.120 142.870 140.120 143.880 ;
        RECT 135.630 142.600 140.120 142.870 ;
        RECT 122.480 141.790 122.740 142.120 ;
        RECT 134.290 141.960 138.780 142.230 ;
        RECT 112.620 141.240 117.110 141.510 ;
        RECT 120.360 141.340 126.160 141.610 ;
        RECT 93.080 140.080 97.030 140.090 ;
        RECT 89.590 139.810 97.030 140.080 ;
        RECT 97.330 140.040 103.130 140.180 ;
        RECT 110.280 140.870 112.280 141.150 ;
        RECT 110.280 140.600 115.770 140.870 ;
        RECT 97.330 139.910 104.580 140.040 ;
        RECT 93.080 139.540 97.030 139.810 ;
        RECT 87.250 139.170 92.740 139.440 ;
        RECT 93.080 139.270 101.830 139.540 ;
        RECT 87.250 138.160 89.250 139.170 ;
        RECT 93.080 138.800 97.030 139.270 ;
        RECT 102.130 138.900 104.580 139.910 ;
        RECT 89.590 138.530 97.030 138.800 ;
        RECT 97.330 138.630 104.580 138.900 ;
        RECT 93.080 138.260 97.030 138.530 ;
        RECT 87.250 137.890 92.740 138.160 ;
        RECT 93.080 138.090 101.830 138.260 ;
        RECT 8.265 137.780 9.275 137.810 ;
        RECT 8.220 136.770 9.320 137.780 ;
        RECT 87.250 136.880 89.250 137.890 ;
        RECT 93.080 137.520 94.080 138.090 ;
        RECT 89.590 137.250 94.080 137.520 ;
        RECT 8.265 136.740 9.275 136.770 ;
        RECT 87.250 136.610 92.740 136.880 ;
        RECT 82.790 134.915 83.860 135.925 ;
        RECT 87.250 135.600 89.250 136.610 ;
        RECT 93.080 136.240 94.080 137.250 ;
        RECT 89.590 135.970 94.080 136.240 ;
        RECT 87.250 135.330 92.740 135.600 ;
        RECT 82.820 133.640 83.830 134.915 ;
        RECT 87.250 134.320 89.250 135.330 ;
        RECT 93.080 134.960 94.080 135.970 ;
        RECT 89.590 134.690 94.080 134.960 ;
        RECT 87.250 134.050 92.740 134.320 ;
        RECT 87.250 133.040 89.250 134.050 ;
        RECT 93.080 133.680 94.080 134.690 ;
        RECT 96.030 137.990 101.830 138.090 ;
        RECT 102.130 138.040 104.580 138.630 ;
        RECT 110.280 139.590 112.280 140.600 ;
        RECT 116.110 140.240 117.110 141.240 ;
        RECT 119.060 140.700 124.860 140.970 ;
        RECT 119.060 140.240 120.060 140.700 ;
        RECT 125.160 140.330 126.160 141.340 ;
        RECT 134.290 141.230 135.290 141.960 ;
        RECT 139.120 141.590 140.120 142.600 ;
        RECT 145.520 142.200 145.720 144.800 ;
        RECT 145.490 141.870 145.750 142.200 ;
        RECT 135.630 141.320 140.120 141.590 ;
        RECT 143.370 141.420 149.170 141.690 ;
        RECT 116.110 140.230 120.060 140.240 ;
        RECT 112.620 139.960 120.060 140.230 ;
        RECT 120.360 140.190 126.160 140.330 ;
        RECT 133.290 140.950 135.290 141.230 ;
        RECT 133.290 140.680 138.780 140.950 ;
        RECT 120.360 140.060 127.610 140.190 ;
        RECT 116.110 139.690 120.060 139.960 ;
        RECT 110.280 139.320 115.770 139.590 ;
        RECT 116.110 139.420 124.860 139.690 ;
        RECT 110.280 138.310 112.280 139.320 ;
        RECT 116.110 138.950 120.060 139.420 ;
        RECT 125.160 139.050 127.610 140.060 ;
        RECT 112.620 138.680 120.060 138.950 ;
        RECT 120.360 138.780 127.610 139.050 ;
        RECT 116.110 138.410 120.060 138.680 ;
        RECT 110.280 138.040 115.770 138.310 ;
        RECT 116.110 138.240 124.860 138.410 ;
        RECT 96.030 136.980 97.030 137.990 ;
        RECT 102.130 137.620 103.130 138.040 ;
        RECT 97.330 137.350 103.130 137.620 ;
        RECT 102.950 137.340 103.130 137.350 ;
        RECT 110.280 137.030 112.280 138.040 ;
        RECT 116.110 137.670 117.110 138.240 ;
        RECT 112.620 137.400 117.110 137.670 ;
        RECT 96.030 136.710 101.830 136.980 ;
        RECT 110.280 136.760 115.770 137.030 ;
        RECT 89.590 133.410 93.420 133.680 ;
        RECT 93.080 133.400 93.420 133.410 ;
        RECT 87.250 131.040 93.700 133.040 ;
        RECT 94.580 130.490 95.780 131.690 ;
        RECT 96.030 128.740 97.030 136.710 ;
        RECT 105.820 135.065 106.890 136.075 ;
        RECT 110.280 135.750 112.280 136.760 ;
        RECT 116.110 136.390 117.110 137.400 ;
        RECT 112.620 136.120 117.110 136.390 ;
        RECT 110.280 135.480 115.770 135.750 ;
        RECT 105.850 133.790 106.860 135.065 ;
        RECT 110.280 134.470 112.280 135.480 ;
        RECT 116.110 135.110 117.110 136.120 ;
        RECT 112.620 134.840 117.110 135.110 ;
        RECT 110.280 134.200 115.770 134.470 ;
        RECT 110.280 133.190 112.280 134.200 ;
        RECT 116.110 133.830 117.110 134.840 ;
        RECT 119.060 138.140 124.860 138.240 ;
        RECT 125.160 138.190 127.610 138.780 ;
        RECT 133.290 139.670 135.290 140.680 ;
        RECT 139.120 140.320 140.120 141.320 ;
        RECT 142.070 140.780 147.870 141.050 ;
        RECT 142.070 140.320 143.070 140.780 ;
        RECT 148.170 140.410 149.170 141.420 ;
        RECT 139.120 140.310 143.070 140.320 ;
        RECT 135.630 140.040 143.070 140.310 ;
        RECT 143.370 140.270 149.170 140.410 ;
        RECT 143.370 140.140 150.620 140.270 ;
        RECT 139.120 139.770 143.070 140.040 ;
        RECT 133.290 139.400 138.780 139.670 ;
        RECT 139.120 139.500 147.870 139.770 ;
        RECT 133.290 138.390 135.290 139.400 ;
        RECT 139.120 139.030 143.070 139.500 ;
        RECT 148.170 139.130 150.620 140.140 ;
        RECT 135.630 138.760 143.070 139.030 ;
        RECT 143.370 138.860 150.620 139.130 ;
        RECT 139.120 138.490 143.070 138.760 ;
        RECT 119.060 137.130 120.060 138.140 ;
        RECT 125.160 137.770 126.160 138.190 ;
        RECT 120.360 137.500 126.160 137.770 ;
        RECT 125.980 137.490 126.160 137.500 ;
        RECT 133.290 138.120 138.780 138.390 ;
        RECT 139.120 138.320 147.870 138.490 ;
        RECT 119.060 136.860 124.860 137.130 ;
        RECT 133.290 137.110 135.290 138.120 ;
        RECT 139.120 137.750 140.120 138.320 ;
        RECT 135.630 137.480 140.120 137.750 ;
        RECT 112.620 133.560 116.450 133.830 ;
        RECT 116.110 133.550 116.450 133.560 ;
        RECT 110.280 131.190 116.730 133.190 ;
        RECT 117.610 130.640 118.810 131.840 ;
        RECT 119.060 128.890 120.060 136.860 ;
        RECT 133.290 136.840 138.780 137.110 ;
        RECT 128.830 135.145 129.900 136.155 ;
        RECT 133.290 135.830 135.290 136.840 ;
        RECT 139.120 136.470 140.120 137.480 ;
        RECT 135.630 136.200 140.120 136.470 ;
        RECT 133.290 135.560 138.780 135.830 ;
        RECT 128.860 133.870 129.870 135.145 ;
        RECT 133.290 134.550 135.290 135.560 ;
        RECT 139.120 135.190 140.120 136.200 ;
        RECT 135.630 134.920 140.120 135.190 ;
        RECT 133.290 134.280 138.780 134.550 ;
        RECT 133.290 133.270 135.290 134.280 ;
        RECT 139.120 133.910 140.120 134.920 ;
        RECT 142.070 138.220 147.870 138.320 ;
        RECT 148.170 138.270 150.620 138.860 ;
        RECT 142.070 137.210 143.070 138.220 ;
        RECT 148.170 137.850 149.170 138.270 ;
        RECT 143.370 137.580 149.170 137.850 ;
        RECT 148.990 137.570 149.170 137.580 ;
        RECT 142.070 136.940 147.870 137.210 ;
        RECT 135.630 133.640 139.460 133.910 ;
        RECT 139.120 133.630 139.460 133.640 ;
        RECT 133.290 131.270 139.740 133.270 ;
        RECT 140.620 130.720 141.820 131.920 ;
        RECT 142.070 129.970 143.070 136.940 ;
        RECT 142.025 128.970 143.115 129.970 ;
        RECT 45.250 29.615 57.010 29.640 ;
        RECT 45.230 28.165 57.010 29.615 ;
        RECT 45.250 28.140 57.010 28.165 ;
        RECT 51.275 18.725 52.600 20.520 ;
        RECT 62.290 20.505 63.610 20.525 ;
        RECT 60.365 19.135 63.635 20.505 ;
        RECT 62.290 19.115 63.610 19.135 ;
        RECT 51.255 17.450 52.620 18.725 ;
        RECT 51.275 17.425 52.600 17.450 ;
        RECT 49.025 12.060 50.475 12.080 ;
        RECT 49.000 10.560 57.140 12.060 ;
        RECT 49.025 10.540 50.475 10.560 ;
      LAYER via2 ;
        RECT 136.060 206.740 137.060 207.740 ;
        RECT 139.760 207.080 140.760 208.080 ;
        RECT 143.440 204.060 144.440 205.060 ;
        RECT 151.540 204.260 152.540 205.260 ;
        RECT 81.850 200.620 82.130 200.900 ;
        RECT 106.590 200.540 106.870 200.820 ;
        RECT 129.840 200.530 130.120 200.810 ;
        RECT 153.470 200.520 153.750 200.800 ;
        RECT 59.625 198.335 60.775 199.485 ;
        RECT 76.150 198.900 76.450 199.190 ;
        RECT 80.200 198.410 81.200 199.410 ;
        RECT 84.365 198.255 85.515 199.405 ;
        RECT 100.890 198.820 101.190 199.110 ;
        RECT 104.940 198.330 105.940 199.330 ;
        RECT 107.615 198.245 108.765 199.395 ;
        RECT 124.140 198.810 124.440 199.100 ;
        RECT 46.620 194.210 47.620 195.210 ;
        RECT 128.190 198.320 129.190 199.320 ;
        RECT 131.245 198.235 132.395 199.385 ;
        RECT 147.770 198.800 148.070 199.090 ;
        RECT 151.820 198.310 152.820 199.310 ;
        RECT 71.350 190.490 73.250 191.330 ;
        RECT 79.350 190.490 81.250 191.330 ;
        RECT 59.540 185.505 60.550 186.515 ;
        RECT 96.090 190.410 97.990 191.250 ;
        RECT 104.090 190.410 105.990 191.250 ;
        RECT 69.110 183.390 70.370 184.830 ;
        RECT 71.400 182.410 72.400 183.410 ;
        RECT 84.280 185.425 85.290 186.435 ;
        RECT 119.340 190.400 121.240 191.240 ;
        RECT 127.340 190.400 129.240 191.240 ;
        RECT 93.850 183.310 95.110 184.750 ;
        RECT 96.140 182.330 97.140 183.330 ;
        RECT 107.530 185.415 108.540 186.425 ;
        RECT 142.970 190.390 144.870 191.230 ;
        RECT 150.970 190.390 152.870 191.230 ;
        RECT 117.100 183.300 118.360 184.740 ;
        RECT 119.390 182.320 120.390 183.320 ;
        RECT 131.160 185.405 132.170 186.415 ;
        RECT 140.730 183.290 141.990 184.730 ;
        RECT 143.020 182.310 144.020 183.310 ;
        RECT 151.860 179.430 152.860 180.430 ;
        RECT 81.740 174.530 82.020 174.810 ;
        RECT 104.920 174.440 105.200 174.720 ;
        RECT 127.820 174.640 128.100 174.920 ;
        RECT 150.920 174.750 151.200 175.030 ;
        RECT 127.820 173.960 128.100 174.240 ;
        RECT 59.515 172.245 60.665 173.395 ;
        RECT 76.040 172.810 76.340 173.100 ;
        RECT 80.090 172.320 81.090 173.320 ;
        RECT 82.695 172.155 83.845 173.305 ;
        RECT 99.220 172.720 99.520 173.010 ;
        RECT 103.270 172.230 104.270 173.230 ;
        RECT 105.595 172.355 106.745 173.505 ;
        RECT 122.120 172.920 122.420 173.210 ;
        RECT 126.170 172.430 127.170 173.430 ;
        RECT 128.695 172.465 129.845 173.615 ;
        RECT 145.220 173.030 145.520 173.320 ;
        RECT 149.270 172.540 150.270 173.540 ;
        RECT 46.990 168.390 47.990 169.390 ;
        RECT 71.240 164.400 73.140 165.240 ;
        RECT 79.240 164.400 81.140 165.240 ;
        RECT 6.745 162.445 7.755 163.455 ;
        RECT 59.430 159.415 60.440 160.425 ;
        RECT 94.420 164.310 96.320 165.150 ;
        RECT 102.420 164.310 104.320 165.150 ;
        RECT 69.000 157.300 70.260 158.740 ;
        RECT 71.290 156.320 72.290 157.320 ;
        RECT 82.610 159.325 83.620 160.335 ;
        RECT 117.320 164.510 119.220 165.350 ;
        RECT 125.320 164.510 127.220 165.350 ;
        RECT 92.180 157.210 93.440 158.650 ;
        RECT 94.470 156.230 95.470 157.230 ;
        RECT 105.510 159.525 106.520 160.535 ;
        RECT 140.420 164.620 142.320 165.460 ;
        RECT 148.420 164.620 150.320 165.460 ;
        RECT 115.080 157.410 116.340 158.850 ;
        RECT 117.370 156.430 118.370 157.430 ;
        RECT 128.610 159.635 129.620 160.645 ;
        RECT 138.180 157.520 139.440 158.960 ;
        RECT 140.470 156.540 141.470 157.540 ;
        RECT 141.820 154.660 142.820 155.660 ;
        RECT 105.130 148.800 105.410 149.080 ;
        RECT 128.160 148.950 128.440 149.230 ;
        RECT 151.170 149.030 151.450 149.310 ;
        RECT 82.905 146.515 84.055 147.665 ;
        RECT 99.430 147.080 99.730 147.370 ;
        RECT 103.480 146.590 104.480 147.590 ;
        RECT 105.935 146.665 107.085 147.815 ;
        RECT 122.460 147.230 122.760 147.520 ;
        RECT 126.510 146.740 127.510 147.740 ;
        RECT 128.945 146.745 130.095 147.895 ;
        RECT 145.470 147.310 145.770 147.600 ;
        RECT 149.520 146.820 150.520 147.820 ;
        RECT 57.170 141.310 58.170 142.310 ;
        RECT 94.630 138.670 96.530 139.510 ;
        RECT 102.630 138.670 104.530 139.510 ;
        RECT 8.265 136.770 9.275 137.780 ;
        RECT 82.820 133.685 83.830 134.695 ;
        RECT 117.660 138.820 119.560 139.660 ;
        RECT 125.660 138.820 127.560 139.660 ;
        RECT 92.390 131.570 93.650 133.010 ;
        RECT 94.680 130.590 95.680 131.590 ;
        RECT 105.850 133.835 106.860 134.845 ;
        RECT 140.670 138.900 142.570 139.740 ;
        RECT 148.670 138.900 150.570 139.740 ;
        RECT 115.420 131.720 116.680 133.160 ;
        RECT 117.710 130.740 118.710 131.740 ;
        RECT 128.860 133.915 129.870 134.925 ;
        RECT 138.430 131.800 139.690 133.240 ;
        RECT 140.720 130.820 141.720 131.820 ;
        RECT 142.070 128.970 143.070 129.970 ;
        RECT 45.275 28.165 46.725 29.615 ;
        RECT 62.290 19.160 63.610 20.480 ;
        RECT 51.300 17.450 52.575 18.725 ;
        RECT 49.025 10.585 50.475 12.035 ;
      LAYER met3 ;
        RECT 139.760 208.105 140.760 209.970 ;
        RECT 136.035 206.715 137.085 207.795 ;
        RECT 139.735 207.055 140.785 208.105 ;
        RECT 143.440 205.085 144.440 206.600 ;
        RECT 151.540 205.285 152.540 207.590 ;
        RECT 143.415 204.035 144.465 205.085 ;
        RECT 151.515 204.235 152.565 205.285 ;
        RECT 81.825 200.595 82.155 200.925 ;
        RECT 59.600 199.505 60.800 199.510 ;
        RECT 59.575 198.315 60.825 199.505 ;
        RECT 76.120 198.870 76.480 199.220 ;
        RECT 59.600 198.310 60.800 198.315 ;
        RECT 46.620 195.235 47.620 196.430 ;
        RECT 76.150 195.660 76.450 198.870 ;
        RECT 80.100 198.310 81.300 199.510 ;
        RECT 81.840 195.660 82.140 200.595 ;
        RECT 106.565 200.515 106.895 200.845 ;
        RECT 84.340 199.425 85.540 199.430 ;
        RECT 84.315 198.235 85.565 199.425 ;
        RECT 100.860 198.790 101.220 199.140 ;
        RECT 84.340 198.230 85.540 198.235 ;
        RECT 76.150 195.360 82.140 195.660 ;
        RECT 100.890 195.580 101.190 198.790 ;
        RECT 104.840 198.230 106.040 199.430 ;
        RECT 106.580 195.580 106.880 200.515 ;
        RECT 129.815 200.505 130.145 200.835 ;
        RECT 107.590 199.415 108.790 199.420 ;
        RECT 107.565 198.225 108.815 199.415 ;
        RECT 124.110 198.780 124.470 199.130 ;
        RECT 107.590 198.220 108.790 198.225 ;
        RECT 100.890 195.280 106.880 195.580 ;
        RECT 124.140 195.570 124.440 198.780 ;
        RECT 128.090 198.220 129.290 199.420 ;
        RECT 129.830 195.570 130.130 200.505 ;
        RECT 153.445 200.495 153.775 200.825 ;
        RECT 131.220 199.405 132.420 199.410 ;
        RECT 131.195 198.215 132.445 199.405 ;
        RECT 147.740 198.770 148.100 199.120 ;
        RECT 131.220 198.210 132.420 198.215 ;
        RECT 124.140 195.270 130.130 195.570 ;
        RECT 147.770 195.560 148.070 198.770 ;
        RECT 151.720 198.210 152.920 199.410 ;
        RECT 153.460 195.560 153.760 200.495 ;
        RECT 147.770 195.260 153.760 195.560 ;
        RECT 46.595 194.185 47.645 195.235 ;
        RECT 71.300 190.460 73.300 191.360 ;
        RECT 79.300 190.460 81.300 191.360 ;
        RECT 4.180 188.235 5.270 189.295 ;
        RECT 59.515 185.480 60.575 186.540 ;
        RECT 59.540 184.245 60.550 185.480 ;
        RECT 79.300 185.310 80.200 190.460 ;
        RECT 96.040 190.380 98.040 191.280 ;
        RECT 104.040 190.380 106.040 191.280 ;
        RECT 84.255 185.400 85.315 186.460 ;
        RECT 69.080 184.410 80.200 185.310 ;
        RECT 69.080 183.360 70.400 184.410 ;
        RECT 84.280 184.165 85.290 185.400 ;
        RECT 104.040 185.230 104.940 190.380 ;
        RECT 119.290 190.370 121.290 191.270 ;
        RECT 127.290 190.370 129.290 191.270 ;
        RECT 107.505 185.390 108.565 186.450 ;
        RECT 93.820 184.330 104.940 185.230 ;
        RECT 71.300 182.310 72.500 183.510 ;
        RECT 93.820 183.280 95.140 184.330 ;
        RECT 107.530 184.155 108.540 185.390 ;
        RECT 127.290 185.220 128.190 190.370 ;
        RECT 142.920 190.360 144.920 191.260 ;
        RECT 150.920 190.360 152.920 191.260 ;
        RECT 131.135 185.380 132.195 186.440 ;
        RECT 117.070 184.320 128.190 185.220 ;
        RECT 96.040 182.230 97.240 183.430 ;
        RECT 117.070 183.270 118.390 184.320 ;
        RECT 131.160 184.145 132.170 185.380 ;
        RECT 150.920 185.210 151.820 190.360 ;
        RECT 140.700 184.310 151.820 185.210 ;
        RECT 119.290 182.220 120.490 183.420 ;
        RECT 140.700 183.260 142.020 184.310 ;
        RECT 142.920 182.210 144.120 183.410 ;
        RECT 127.770 179.090 128.150 179.410 ;
        RECT 151.835 179.405 152.885 180.455 ;
        RECT 81.720 176.830 82.040 177.210 ;
        RECT 81.730 174.835 82.030 176.830 ;
        RECT 104.900 176.280 105.220 176.660 ;
        RECT 81.715 174.505 82.045 174.835 ;
        RECT 104.910 174.745 105.210 176.280 ;
        RECT 127.810 174.945 128.110 179.090 ;
        RECT 150.870 178.240 151.250 178.560 ;
        RECT 151.860 178.240 152.860 179.405 ;
        RECT 150.910 175.055 151.210 178.240 ;
        RECT 59.490 173.415 60.690 173.420 ;
        RECT 59.465 172.225 60.715 173.415 ;
        RECT 76.010 172.780 76.370 173.130 ;
        RECT 59.490 172.220 60.690 172.225 ;
        RECT 76.040 169.570 76.340 172.780 ;
        RECT 79.990 172.220 81.190 173.420 ;
        RECT 81.730 169.570 82.030 174.505 ;
        RECT 104.895 174.415 105.225 174.745 ;
        RECT 127.795 174.615 128.125 174.945 ;
        RECT 150.895 174.725 151.225 175.055 ;
        RECT 82.670 173.325 83.870 173.330 ;
        RECT 82.645 172.135 83.895 173.325 ;
        RECT 99.190 172.690 99.550 173.040 ;
        RECT 82.670 172.130 83.870 172.135 ;
        RECT 46.965 168.365 48.015 169.445 ;
        RECT 76.040 169.270 82.030 169.570 ;
        RECT 99.220 169.480 99.520 172.690 ;
        RECT 103.170 172.130 104.370 173.330 ;
        RECT 104.910 169.480 105.210 174.415 ;
        RECT 127.810 174.265 128.110 174.615 ;
        RECT 127.795 173.935 128.125 174.265 ;
        RECT 105.570 173.525 106.770 173.530 ;
        RECT 105.545 172.335 106.795 173.525 ;
        RECT 122.090 172.890 122.450 173.240 ;
        RECT 105.570 172.330 106.770 172.335 ;
        RECT 99.220 169.180 105.210 169.480 ;
        RECT 122.120 169.680 122.420 172.890 ;
        RECT 126.070 172.330 127.270 173.530 ;
        RECT 127.810 169.680 128.110 173.935 ;
        RECT 128.670 173.635 129.870 173.640 ;
        RECT 128.645 172.445 129.895 173.635 ;
        RECT 145.190 173.000 145.550 173.350 ;
        RECT 128.670 172.440 129.870 172.445 ;
        RECT 122.120 169.380 128.110 169.680 ;
        RECT 145.220 169.790 145.520 173.000 ;
        RECT 149.170 172.440 150.370 173.640 ;
        RECT 150.910 169.790 151.210 174.725 ;
        RECT 145.220 169.490 151.210 169.790 ;
        RECT 71.190 164.370 73.190 165.270 ;
        RECT 79.190 164.370 81.190 165.270 ;
        RECT 6.720 163.455 7.780 163.480 ;
        RECT 4.975 162.445 7.780 163.455 ;
        RECT 6.720 162.420 7.780 162.445 ;
        RECT 59.405 159.390 60.465 160.450 ;
        RECT 59.430 158.155 60.440 159.390 ;
        RECT 79.190 159.220 80.090 164.370 ;
        RECT 94.370 164.280 96.370 165.180 ;
        RECT 102.370 164.280 104.370 165.180 ;
        RECT 117.270 164.480 119.270 165.380 ;
        RECT 125.270 164.480 127.270 165.380 ;
        RECT 140.370 164.590 142.370 165.490 ;
        RECT 148.370 164.590 150.370 165.490 ;
        RECT 82.585 159.300 83.645 160.360 ;
        RECT 68.970 158.320 80.090 159.220 ;
        RECT 68.970 157.270 70.290 158.320 ;
        RECT 82.610 158.065 83.620 159.300 ;
        RECT 102.370 159.130 103.270 164.280 ;
        RECT 105.485 159.500 106.545 160.560 ;
        RECT 92.150 158.230 103.270 159.130 ;
        RECT 105.510 158.265 106.520 159.500 ;
        RECT 125.270 159.330 126.170 164.480 ;
        RECT 128.585 159.610 129.645 160.670 ;
        RECT 115.050 158.430 126.170 159.330 ;
        RECT 71.190 156.220 72.390 157.420 ;
        RECT 92.150 157.180 93.470 158.230 ;
        RECT 115.050 157.380 116.370 158.430 ;
        RECT 128.610 158.375 129.620 159.610 ;
        RECT 148.370 159.440 149.270 164.590 ;
        RECT 138.150 158.540 149.270 159.440 ;
        RECT 94.370 156.130 95.570 157.330 ;
        RECT 117.270 156.330 118.470 157.530 ;
        RECT 138.150 157.490 139.470 158.540 ;
        RECT 140.370 156.440 141.570 157.640 ;
        RECT 141.795 155.660 142.845 155.685 ;
        RECT 141.795 154.660 149.940 155.660 ;
        RECT 141.795 154.635 142.845 154.660 ;
        RECT 128.140 152.490 128.460 152.870 ;
        RECT 105.110 150.650 105.430 151.030 ;
        RECT 105.120 149.105 105.420 150.650 ;
        RECT 128.150 149.255 128.450 152.490 ;
        RECT 151.150 151.450 151.470 151.830 ;
        RECT 151.160 149.335 151.460 151.450 ;
        RECT 105.105 148.775 105.435 149.105 ;
        RECT 128.135 148.925 128.465 149.255 ;
        RECT 151.145 149.005 151.475 149.335 ;
        RECT 82.880 147.685 84.080 147.690 ;
        RECT 82.855 146.495 84.105 147.685 ;
        RECT 99.400 147.050 99.760 147.400 ;
        RECT 82.880 146.490 84.080 146.495 ;
        RECT 99.430 143.840 99.730 147.050 ;
        RECT 103.380 146.490 104.580 147.690 ;
        RECT 105.120 143.840 105.420 148.775 ;
        RECT 105.910 147.835 107.110 147.840 ;
        RECT 105.885 146.645 107.135 147.835 ;
        RECT 122.430 147.200 122.790 147.550 ;
        RECT 105.910 146.640 107.110 146.645 ;
        RECT 99.430 143.540 105.420 143.840 ;
        RECT 122.460 143.990 122.760 147.200 ;
        RECT 126.410 146.640 127.610 147.840 ;
        RECT 128.150 143.990 128.450 148.925 ;
        RECT 128.920 147.915 130.120 147.920 ;
        RECT 128.895 146.725 130.145 147.915 ;
        RECT 145.440 147.280 145.800 147.630 ;
        RECT 128.920 146.720 130.120 146.725 ;
        RECT 122.460 143.690 128.450 143.990 ;
        RECT 145.470 144.070 145.770 147.280 ;
        RECT 149.420 146.720 150.620 147.920 ;
        RECT 151.160 144.070 151.460 149.005 ;
        RECT 145.470 143.770 151.460 144.070 ;
        RECT 57.115 141.285 58.195 142.335 ;
        RECT 94.580 138.640 96.580 139.540 ;
        RECT 102.580 138.640 104.580 139.540 ;
        RECT 117.610 138.790 119.610 139.690 ;
        RECT 125.610 138.790 127.610 139.690 ;
        RECT 140.620 138.870 142.620 139.770 ;
        RECT 148.620 138.870 150.620 139.770 ;
        RECT 8.240 137.780 9.300 137.805 ;
        RECT 5.815 136.770 9.300 137.780 ;
        RECT 8.240 136.745 9.300 136.770 ;
        RECT 82.795 133.660 83.855 134.720 ;
        RECT 82.820 132.425 83.830 133.660 ;
        RECT 102.580 133.490 103.480 138.640 ;
        RECT 105.825 133.810 106.885 134.870 ;
        RECT 92.360 132.590 103.480 133.490 ;
        RECT 92.360 131.540 93.680 132.590 ;
        RECT 105.850 132.575 106.860 133.810 ;
        RECT 125.610 133.640 126.510 138.790 ;
        RECT 128.835 133.890 129.895 134.950 ;
        RECT 115.390 132.740 126.510 133.640 ;
        RECT 115.390 131.690 116.710 132.740 ;
        RECT 128.860 132.655 129.870 133.890 ;
        RECT 148.620 133.720 149.520 138.870 ;
        RECT 138.400 132.820 149.520 133.720 ;
        RECT 94.580 130.490 95.780 131.690 ;
        RECT 117.610 130.640 118.810 131.840 ;
        RECT 138.400 131.770 139.720 132.820 ;
        RECT 140.620 130.720 141.820 131.920 ;
        RECT 142.045 129.970 143.095 129.995 ;
        RECT 147.160 129.970 148.160 130.000 ;
        RECT 142.045 128.970 148.160 129.970 ;
        RECT 142.045 128.945 143.095 128.970 ;
        RECT 147.160 128.940 148.160 128.970 ;
        RECT 45.255 29.640 46.745 29.665 ;
        RECT 45.250 28.140 46.750 29.640 ;
        RECT 45.255 28.115 46.745 28.140 ;
        RECT 62.265 20.500 63.635 20.505 ;
        RECT 62.240 19.140 63.660 20.500 ;
        RECT 62.265 19.135 63.635 19.140 ;
        RECT 51.275 18.745 52.600 18.750 ;
        RECT 51.250 17.430 52.625 18.745 ;
        RECT 51.275 17.425 52.600 17.430 ;
        RECT 49.005 12.060 50.495 12.085 ;
        RECT 49.000 10.560 50.500 12.060 ;
        RECT 49.005 10.535 50.495 10.560 ;
      LAYER via3 ;
        RECT 139.760 208.940 140.760 209.940 ;
        RECT 136.035 206.765 137.085 207.765 ;
        RECT 143.440 205.570 144.440 206.570 ;
        RECT 151.540 206.560 152.540 207.560 ;
        RECT 59.605 198.315 60.795 199.505 ;
        RECT 46.620 195.400 47.620 196.400 ;
        RECT 80.200 198.410 81.200 199.410 ;
        RECT 84.345 198.235 85.535 199.425 ;
        RECT 104.940 198.330 105.940 199.330 ;
        RECT 107.595 198.225 108.785 199.415 ;
        RECT 128.190 198.320 129.190 199.320 ;
        RECT 131.225 198.215 132.415 199.405 ;
        RECT 151.820 198.310 152.820 199.310 ;
        RECT 71.330 190.490 73.270 191.330 ;
        RECT 79.330 190.490 81.270 191.330 ;
        RECT 4.210 188.235 5.220 189.295 ;
        RECT 96.070 190.410 98.010 191.250 ;
        RECT 104.070 190.410 106.010 191.250 ;
        RECT 119.320 190.400 121.260 191.240 ;
        RECT 59.540 184.275 60.550 185.285 ;
        RECT 127.320 190.400 129.260 191.240 ;
        RECT 142.950 190.390 144.890 191.230 ;
        RECT 84.280 184.195 85.290 185.205 ;
        RECT 150.950 190.390 152.890 191.230 ;
        RECT 71.400 182.410 72.400 183.410 ;
        RECT 107.530 184.185 108.540 185.195 ;
        RECT 96.140 182.330 97.140 183.330 ;
        RECT 131.160 184.175 132.170 185.185 ;
        RECT 119.390 182.320 120.390 183.320 ;
        RECT 143.020 182.310 144.020 183.310 ;
        RECT 127.800 179.090 128.120 179.410 ;
        RECT 81.720 176.860 82.040 177.180 ;
        RECT 104.900 176.310 105.220 176.630 ;
        RECT 150.900 178.240 151.220 178.560 ;
        RECT 151.860 178.270 152.860 179.270 ;
        RECT 59.495 172.225 60.685 173.415 ;
        RECT 80.090 172.320 81.090 173.320 ;
        RECT 82.675 172.135 83.865 173.325 ;
        RECT 46.965 168.415 48.015 169.415 ;
        RECT 103.270 172.230 104.270 173.230 ;
        RECT 105.575 172.335 106.765 173.525 ;
        RECT 126.170 172.430 127.170 173.430 ;
        RECT 128.675 172.445 129.865 173.635 ;
        RECT 149.270 172.540 150.270 173.540 ;
        RECT 71.220 164.400 73.160 165.240 ;
        RECT 79.220 164.400 81.160 165.240 ;
        RECT 5.005 162.445 6.015 163.455 ;
        RECT 94.400 164.310 96.340 165.150 ;
        RECT 102.400 164.310 104.340 165.150 ;
        RECT 117.300 164.510 119.240 165.350 ;
        RECT 125.300 164.510 127.240 165.350 ;
        RECT 140.400 164.620 142.340 165.460 ;
        RECT 148.400 164.620 150.340 165.460 ;
        RECT 59.430 158.185 60.440 159.195 ;
        RECT 82.610 158.095 83.620 159.105 ;
        RECT 105.510 158.295 106.520 159.305 ;
        RECT 71.290 156.320 72.290 157.320 ;
        RECT 128.610 158.405 129.620 159.415 ;
        RECT 94.470 156.230 95.470 157.230 ;
        RECT 117.370 156.430 118.370 157.430 ;
        RECT 140.470 156.540 141.470 157.540 ;
        RECT 148.910 154.660 149.910 155.660 ;
        RECT 128.140 152.520 128.460 152.840 ;
        RECT 105.110 150.680 105.430 151.000 ;
        RECT 151.150 151.480 151.470 151.800 ;
        RECT 82.885 146.495 84.075 147.685 ;
        RECT 103.480 146.590 104.480 147.590 ;
        RECT 105.915 146.645 107.105 147.835 ;
        RECT 126.510 146.740 127.510 147.740 ;
        RECT 128.925 146.725 130.115 147.915 ;
        RECT 149.520 146.820 150.520 147.820 ;
        RECT 57.145 141.285 58.145 142.335 ;
        RECT 94.610 138.670 96.550 139.510 ;
        RECT 102.610 138.670 104.550 139.510 ;
        RECT 117.640 138.820 119.580 139.660 ;
        RECT 125.640 138.820 127.580 139.660 ;
        RECT 140.650 138.900 142.590 139.740 ;
        RECT 148.650 138.900 150.590 139.740 ;
        RECT 5.845 136.770 6.855 137.780 ;
        RECT 82.820 132.455 83.830 133.465 ;
        RECT 105.850 132.605 106.860 133.615 ;
        RECT 128.860 132.685 129.870 133.695 ;
        RECT 94.680 130.590 95.680 131.590 ;
        RECT 117.710 130.740 118.710 131.740 ;
        RECT 140.720 130.820 141.720 131.820 ;
        RECT 147.160 128.970 148.160 129.970 ;
        RECT 45.255 28.145 46.745 29.635 ;
        RECT 62.270 19.140 63.630 20.500 ;
        RECT 51.280 17.430 52.595 18.745 ;
        RECT 49.005 10.565 50.495 12.055 ;
      LAYER met4 ;
        RECT 110.690 224.760 110.710 225.330 ;
        RECT 114.360 224.760 114.390 225.550 ;
        RECT 136.060 224.760 136.470 225.760 ;
        RECT 136.770 224.760 137.060 225.760 ;
        RECT 139.755 225.150 140.150 225.760 ;
        RECT 3.990 223.390 4.290 224.760 ;
        RECT 7.670 223.390 7.970 224.760 ;
        RECT 11.350 223.390 11.650 224.760 ;
        RECT 15.030 223.390 15.330 224.760 ;
        RECT 18.710 223.390 19.010 224.760 ;
        RECT 22.390 223.390 22.690 224.760 ;
        RECT 26.070 223.390 26.370 224.760 ;
        RECT 29.750 223.390 30.050 224.760 ;
        RECT 33.430 223.390 33.730 224.760 ;
        RECT 37.110 223.390 37.410 224.760 ;
        RECT 40.790 223.390 41.090 224.760 ;
        RECT 44.470 223.390 44.770 224.760 ;
        RECT 48.150 223.390 48.450 224.760 ;
        RECT 51.830 223.390 52.130 224.760 ;
        RECT 55.510 223.390 55.810 224.760 ;
        RECT 59.190 223.390 59.490 224.760 ;
        RECT 62.870 223.390 63.170 224.760 ;
        RECT 66.550 223.390 66.850 224.760 ;
        RECT 70.230 223.390 70.530 224.760 ;
        RECT 73.910 223.390 74.210 224.760 ;
        RECT 77.590 223.390 77.890 224.760 ;
        RECT 81.270 223.390 81.570 224.760 ;
        RECT 84.950 223.390 85.250 224.760 ;
        RECT 88.630 223.390 88.930 224.760 ;
        RECT 3.385 222.320 89.730 223.390 ;
        RECT 49.000 220.760 50.500 222.320 ;
        RECT 59.170 222.300 59.490 222.320 ;
        RECT 110.690 209.660 110.990 224.760 ;
        RECT 97.860 209.360 110.990 209.660 ;
        RECT 97.860 208.190 98.160 209.360 ;
        RECT 114.360 208.900 114.660 224.760 ;
        RECT 74.480 207.890 98.160 208.190 ;
        RECT 98.690 208.600 114.660 208.900 ;
        RECT 46.615 196.400 47.625 196.405 ;
        RECT 46.615 195.400 49.000 196.400 ;
        RECT 46.615 195.395 47.625 195.400 ;
        RECT 50.500 192.800 50.790 193.800 ;
        RECT 4.205 189.270 5.225 189.300 ;
        RECT 2.500 188.260 5.225 189.270 ;
        RECT 4.205 188.230 5.225 188.260 ;
        RECT 46.960 169.415 48.020 169.420 ;
        RECT 46.960 168.415 49.000 169.415 ;
        RECT 46.960 168.410 48.020 168.415 ;
        RECT 50.500 167.030 50.520 168.030 ;
        RECT 5.000 163.455 6.020 163.460 ;
        RECT 2.500 162.445 6.020 163.455 ;
        RECT 5.000 162.440 6.020 162.445 ;
        RECT 52.900 150.960 53.200 206.870 ;
        RECT 74.480 205.540 74.780 207.890 ;
        RECT 98.690 207.410 98.990 208.600 ;
        RECT 118.070 208.180 118.370 224.760 ;
        RECT 121.750 209.160 122.050 224.760 ;
        RECT 54.010 205.240 74.780 205.540 ;
        RECT 75.460 207.110 98.990 207.410 ;
        RECT 99.430 207.880 118.370 208.180 ;
        RECT 121.380 208.860 122.050 209.160 ;
        RECT 54.010 151.910 54.310 205.240 ;
        RECT 75.460 204.570 75.760 207.110 ;
        RECT 99.430 206.430 99.730 207.880 ;
        RECT 121.380 207.480 121.680 208.860 ;
        RECT 125.430 208.480 125.730 224.760 ;
        RECT 55.080 204.270 75.760 204.570 ;
        RECT 76.510 206.130 99.730 206.430 ;
        RECT 100.150 207.180 121.680 207.480 ;
        RECT 122.180 208.180 125.730 208.480 ;
        RECT 55.080 152.840 55.380 204.270 ;
        RECT 59.170 203.440 59.490 203.450 ;
        RECT 55.930 203.360 59.490 203.440 ;
        RECT 76.510 203.360 76.810 206.130 ;
        RECT 100.150 205.750 100.450 207.180 ;
        RECT 122.180 206.770 122.480 208.180 ;
        RECT 129.110 207.680 129.410 224.760 ;
        RECT 55.930 203.120 76.810 203.360 ;
        RECT 55.930 153.710 56.250 203.120 ;
        RECT 59.220 203.060 76.810 203.120 ;
        RECT 77.180 205.450 100.450 205.750 ;
        RECT 100.860 206.470 122.480 206.770 ;
        RECT 122.850 207.380 129.410 207.680 ;
        RECT 77.180 202.710 77.480 205.450 ;
        RECT 100.860 205.050 101.160 206.470 ;
        RECT 122.850 205.990 123.150 207.380 ;
        RECT 132.790 206.970 133.090 224.760 ;
        RECT 136.060 207.770 137.060 224.760 ;
        RECT 139.760 224.760 140.150 225.150 ;
        RECT 140.450 224.760 140.760 225.760 ;
        RECT 139.760 209.945 140.760 224.760 ;
        RECT 143.440 224.760 143.830 225.760 ;
        RECT 144.130 224.760 144.440 225.760 ;
        RECT 139.755 208.935 140.765 209.945 ;
        RECT 56.610 202.410 77.480 202.710 ;
        RECT 77.830 204.750 101.160 205.050 ;
        RECT 101.520 205.690 123.150 205.990 ;
        RECT 123.560 206.670 133.090 206.970 ;
        RECT 136.030 206.760 137.090 207.770 ;
        RECT 56.610 178.070 56.910 202.410 ;
        RECT 77.830 202.030 78.130 204.750 ;
        RECT 101.520 204.270 101.820 205.690 ;
        RECT 123.560 205.370 123.860 206.670 ;
        RECT 143.440 206.575 144.440 224.760 ;
        RECT 147.110 224.760 147.510 225.760 ;
        RECT 147.810 224.760 148.110 225.760 ;
        RECT 147.110 207.560 148.110 224.760 ;
        RECT 151.535 207.560 152.545 207.565 ;
        RECT 143.435 205.565 144.445 206.575 ;
        RECT 147.110 206.560 152.545 207.560 ;
        RECT 151.535 206.555 152.545 206.560 ;
        RECT 57.270 201.730 78.130 202.030 ;
        RECT 78.640 203.970 101.820 204.270 ;
        RECT 102.160 205.070 123.860 205.370 ;
        RECT 57.270 178.670 57.570 201.730 ;
        RECT 78.640 201.230 78.940 203.970 ;
        RECT 102.160 203.500 102.460 205.070 ;
        RECT 57.920 200.930 78.940 201.230 ;
        RECT 79.300 203.200 102.460 203.500 ;
        RECT 57.920 179.410 58.220 200.930 ;
        RECT 79.300 200.490 79.600 203.200 ;
        RECT 58.630 200.190 79.600 200.490 ;
        RECT 58.630 180.030 58.930 200.190 ;
        RECT 59.540 199.430 81.300 199.510 ;
        RECT 59.540 199.420 106.040 199.430 ;
        RECT 59.540 199.410 132.490 199.420 ;
        RECT 59.540 198.310 152.920 199.410 ;
        RECT 80.150 198.230 152.920 198.310 ;
        RECT 104.720 198.220 152.920 198.230 ;
        RECT 131.160 198.210 152.920 198.220 ;
        RECT 71.300 190.460 73.300 191.360 ;
        RECT 79.300 190.460 81.300 191.360 ;
        RECT 96.040 190.380 98.040 191.280 ;
        RECT 104.040 190.380 106.040 191.280 ;
        RECT 119.290 190.370 121.290 191.270 ;
        RECT 127.290 190.370 129.290 191.270 ;
        RECT 142.920 190.360 144.920 191.260 ;
        RECT 150.920 190.360 152.920 191.260 ;
        RECT 59.535 184.270 60.555 185.290 ;
        RECT 59.540 183.510 60.550 184.270 ;
        RECT 84.275 184.190 85.295 185.210 ;
        RECT 59.540 183.430 81.300 183.510 ;
        RECT 84.280 183.430 85.290 184.190 ;
        RECT 107.525 184.180 108.545 185.200 ;
        RECT 59.540 183.420 106.040 183.430 ;
        RECT 107.530 183.420 108.540 184.180 ;
        RECT 131.155 184.170 132.175 185.190 ;
        RECT 131.160 183.420 132.170 184.170 ;
        RECT 59.540 183.410 133.400 183.420 ;
        RECT 59.540 182.310 152.920 183.410 ;
        RECT 76.130 182.230 152.920 182.310 ;
        RECT 101.070 182.220 152.920 182.230 ;
        RECT 131.160 182.210 152.920 182.220 ;
        RECT 58.630 179.730 151.210 180.030 ;
        RECT 57.920 179.400 126.030 179.410 ;
        RECT 127.795 179.400 128.125 179.415 ;
        RECT 57.920 179.110 128.125 179.400 ;
        RECT 125.680 179.100 128.125 179.110 ;
        RECT 127.795 179.085 128.125 179.100 ;
        RECT 57.270 178.370 105.210 178.670 ;
        RECT 150.910 178.565 151.210 179.730 ;
        RECT 56.610 178.060 80.480 178.070 ;
        RECT 56.610 177.770 82.030 178.060 ;
        RECT 80.230 177.760 82.030 177.770 ;
        RECT 81.730 177.185 82.030 177.760 ;
        RECT 81.715 176.855 82.045 177.185 ;
        RECT 104.910 176.635 105.210 178.370 ;
        RECT 150.895 178.235 151.225 178.565 ;
        RECT 151.855 178.265 152.865 179.275 ;
        RECT 104.895 176.305 105.225 176.635 ;
        RECT 126.160 173.530 150.370 173.640 ;
        RECT 59.430 173.330 81.190 173.420 ;
        RECT 103.230 173.330 150.370 173.530 ;
        RECT 59.430 172.440 150.370 173.330 ;
        RECT 59.430 172.330 127.270 172.440 ;
        RECT 59.430 172.220 104.370 172.330 ;
        RECT 80.040 172.130 104.370 172.220 ;
        RECT 71.190 164.370 73.190 165.270 ;
        RECT 79.190 164.370 81.190 165.270 ;
        RECT 94.370 164.280 96.370 165.180 ;
        RECT 102.370 164.280 104.370 165.180 ;
        RECT 117.270 164.480 119.270 165.380 ;
        RECT 125.270 164.480 127.270 165.380 ;
        RECT 140.370 164.590 142.370 165.490 ;
        RECT 148.370 164.590 150.370 165.490 ;
        RECT 59.425 158.180 60.445 159.200 ;
        RECT 59.430 157.420 60.440 158.180 ;
        RECT 82.605 158.090 83.625 159.110 ;
        RECT 105.505 158.290 106.525 159.310 ;
        RECT 128.605 158.400 129.625 159.420 ;
        RECT 59.430 157.330 81.190 157.420 ;
        RECT 82.610 157.330 83.620 158.090 ;
        RECT 105.510 157.530 106.520 158.290 ;
        RECT 128.610 157.640 129.620 158.400 ;
        RECT 122.120 157.530 150.370 157.640 ;
        RECT 101.060 157.330 150.370 157.530 ;
        RECT 59.430 156.440 150.370 157.330 ;
        RECT 59.430 156.330 127.270 156.440 ;
        RECT 59.430 156.220 104.370 156.330 ;
        RECT 76.290 156.130 104.370 156.220 ;
        RECT 148.905 155.660 149.915 155.665 ;
        RECT 151.860 155.660 152.860 178.265 ;
        RECT 148.905 154.660 152.860 155.660 ;
        RECT 148.905 154.655 149.915 154.660 ;
        RECT 55.930 153.390 151.460 153.710 ;
        RECT 55.080 152.830 127.700 152.840 ;
        RECT 128.135 152.830 128.465 152.845 ;
        RECT 55.080 152.540 128.465 152.830 ;
        RECT 127.350 152.530 128.465 152.540 ;
        RECT 128.135 152.515 128.465 152.530 ;
        RECT 105.120 151.910 105.420 151.940 ;
        RECT 54.010 151.610 105.420 151.910 ;
        RECT 151.160 151.805 151.460 153.390 ;
        RECT 105.120 151.005 105.420 151.610 ;
        RECT 151.145 151.475 151.475 151.805 ;
        RECT 52.900 150.660 82.020 150.960 ;
        RECT 105.105 150.675 105.435 151.005 ;
        RECT 126.390 147.840 150.620 147.920 ;
        RECT 103.390 147.690 150.620 147.840 ;
        RECT 82.820 146.720 150.620 147.690 ;
        RECT 82.820 146.640 127.610 146.720 ;
        RECT 82.820 146.490 104.580 146.640 ;
        RECT 57.140 142.310 58.150 142.340 ;
        RECT 50.500 141.310 58.150 142.310 ;
        RECT 57.140 141.280 58.150 141.310 ;
        RECT 94.580 138.640 96.580 139.540 ;
        RECT 102.580 138.640 104.580 139.540 ;
        RECT 117.610 138.790 119.610 139.690 ;
        RECT 125.610 138.790 127.610 139.690 ;
        RECT 140.620 138.870 142.620 139.770 ;
        RECT 148.620 138.870 150.620 139.770 ;
        RECT 5.840 137.780 6.860 137.785 ;
        RECT 2.500 136.770 6.860 137.780 ;
        RECT 5.840 136.765 6.860 136.770 ;
        RECT 82.815 132.450 83.835 133.470 ;
        RECT 105.845 132.600 106.865 133.620 ;
        RECT 128.855 132.680 129.875 133.700 ;
        RECT 82.820 131.690 83.830 132.450 ;
        RECT 105.850 131.840 106.860 132.600 ;
        RECT 128.860 131.920 129.870 132.680 ;
        RECT 122.440 131.840 150.620 131.920 ;
        RECT 98.260 131.690 150.620 131.840 ;
        RECT 82.820 130.720 150.620 131.690 ;
        RECT 82.820 130.640 127.610 130.720 ;
        RECT 82.820 130.490 104.580 130.640 ;
        RECT 147.155 129.970 148.165 129.975 ;
        RECT 151.860 129.970 152.860 154.660 ;
        RECT 147.155 128.970 152.860 129.970 ;
        RECT 147.155 128.965 148.165 128.970 ;
        RECT 2.500 36.100 43.370 37.600 ;
        RECT 41.870 29.640 43.370 36.100 ;
        RECT 41.870 28.140 46.750 29.640 ;
        RECT 49.000 2.310 50.500 5.000 ;
        RECT 51.275 1.365 52.600 18.750 ;
        RECT 45.800 1.000 52.600 1.365 ;
        RECT 45.800 0.600 46.160 1.000 ;
        RECT 45.790 0.000 46.160 0.600 ;
        RECT 46.760 0.000 52.600 1.000 ;
        RECT 62.265 1.385 63.635 20.505 ;
        RECT 151.860 3.220 152.860 128.970 ;
        RECT 151.860 2.220 157.060 3.220 ;
        RECT 62.265 1.000 69.225 1.385 ;
        RECT 156.060 1.140 157.060 2.220 ;
        RECT 62.265 0.600 68.240 1.000 ;
        RECT 62.260 0.000 68.240 0.600 ;
        RECT 68.840 0.600 69.225 1.000 ;
        RECT 156.000 1.000 157.160 1.140 ;
        RECT 68.840 0.000 69.230 0.600 ;
        RECT 156.000 0.000 156.560 1.000 ;
  END
END tt_um_JamesTimothyMeech_inverter
END LIBRARY

