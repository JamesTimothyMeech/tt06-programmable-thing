** sch_path: /home/james/Desktop/TinyTapeout/TinyTapeoutAnalog/tt_asw_1v8/xschem/analog_mux.sch
.subckt analog_mux VPWR ctrl mod bus VGND
*.PININFO VPWR:B VGND:B mod:B bus:B ctrl:I
XM4 tgon tgon_n VGND VGND sky130_fd_pr__nfet_01v8 L=0.15 W=1.5 nf=1 m=1
XM3 tgon tgon_n VPWR VPWR sky130_fd_pr__pfet_01v8 L=0.15 W=3 nf=2 m=1
XM2 tgon_n ctrl VGND VGND sky130_fd_pr__nfet_01v8 L=0.15 W=1.5 nf=1 m=1
XM1 tgon_n ctrl VPWR VPWR sky130_fd_pr__pfet_01v8 L=0.15 W=3 nf=2 m=1
XM6 bus tgon mod VGND sky130_fd_pr__nfet_01v8_lvt L=0.35 W=31.5 nf=7 m=1
XM5 bus tgon_n mod VPWR sky130_fd_pr__pfet_01v8_lvt L=0.35 W=94.5 nf=21 m=1
XR1 VGND mod VGND sky130_fd_pr__res_xhigh_po_0p35 L=10 mult=1 m=1
.ends
.end
