magic
tech sky130A
magscale 1 2
timestamp 1713457832
<< metal1 >>
rect 30308 40674 30508 40680
rect 30308 40042 30508 40474
rect 25820 38560 25826 38760
rect 26026 38560 26416 38760
rect 1365 37652 1371 37854
rect 1573 37652 26434 37854
rect 28588 36104 30372 36304
rect 30572 36104 30578 36304
rect 11096 5928 11396 6474
rect 11096 5622 11396 5628
rect 12079 4101 12353 4107
rect 10249 3833 10255 4098
rect 10520 3833 10870 4098
rect 12079 3821 12353 3827
rect 11122 2412 11422 2418
rect 11122 1730 11422 2112
<< via1 >>
rect 30308 40474 30508 40674
rect 25826 38560 26026 38760
rect 1371 37652 1573 37854
rect 30372 36104 30572 36304
rect 11096 5628 11396 5928
rect 10255 3833 10520 4098
rect 12079 3827 12353 4101
rect 11122 2112 11422 2412
<< metal2 >>
rect 30308 41052 30508 41061
rect 30308 40674 30508 40852
rect 30302 40474 30308 40674
rect 30508 40474 30514 40674
rect 25826 38760 26026 38766
rect 25599 38560 25608 38760
rect 25808 38560 25826 38760
rect 25826 38554 26026 38560
rect 847 37854 1049 37863
rect 1371 37854 1573 37860
rect 1049 37652 1371 37854
rect 847 37643 1049 37652
rect 1371 37646 1573 37652
rect 30372 36304 30572 36310
rect 30372 36086 30572 36104
rect 30372 35877 30572 35886
rect 9050 5923 11096 5928
rect 9046 5633 9055 5923
rect 9345 5633 11096 5923
rect 9050 5628 11096 5633
rect 11396 5628 11402 5928
rect 10255 4098 10520 4104
rect 12458 4101 12722 4105
rect 10255 3745 10520 3833
rect 12073 3827 12079 4101
rect 12353 4096 12727 4101
rect 12353 3832 12458 4096
rect 12722 3832 12727 4096
rect 12353 3827 12727 3832
rect 12458 3823 12722 3827
rect 10251 3490 10260 3745
rect 10515 3490 10524 3745
rect 10255 3485 10520 3490
rect 9805 2412 10095 2416
rect 9800 2407 11122 2412
rect 9800 2117 9805 2407
rect 10095 2117 11122 2407
rect 9800 2112 11122 2117
rect 11422 2112 11428 2412
rect 9805 2108 10095 2112
<< via2 >>
rect 30308 40852 30508 41052
rect 25608 38560 25808 38760
rect 847 37652 1049 37854
rect 30372 35886 30572 36086
rect 9055 5633 9345 5923
rect 12458 3832 12722 4096
rect 10260 3490 10515 3745
rect 9805 2117 10095 2407
<< metal3 >>
rect 30308 41512 30508 41518
rect 30308 41057 30508 41312
rect 30303 41052 30513 41057
rect 30303 40852 30308 41052
rect 30508 40852 30513 41052
rect 30303 40847 30513 40852
rect 25603 38760 25813 38765
rect 25376 38560 25382 38760
rect 25582 38560 25608 38760
rect 25808 38560 25813 38760
rect 25603 38555 25813 38560
rect 836 37647 842 37859
rect 1044 37854 1054 37859
rect 1049 37652 1054 37854
rect 1044 37647 1054 37652
rect 30367 36086 30577 36091
rect 30367 35886 30372 36086
rect 30572 35886 30577 36086
rect 30367 35881 30577 35886
rect 30372 35854 30572 35881
rect 30372 35648 30572 35654
rect 9051 5928 9349 5933
rect 9050 5927 9350 5928
rect 9050 5629 9051 5927
rect 9349 5629 9350 5927
rect 9050 5628 9350 5629
rect 9051 5623 9349 5628
rect 12453 4100 12727 4101
rect 12448 3828 12454 4100
rect 12726 3828 12732 4100
rect 12453 3827 12727 3828
rect 10255 3749 10520 3750
rect 10250 3486 10256 3749
rect 10519 3486 10525 3749
rect 10255 3485 10520 3486
rect 9801 2412 10099 2417
rect 9800 2411 10100 2412
rect 9800 2113 9801 2411
rect 10099 2113 10100 2411
rect 9800 2112 10100 2113
rect 9801 2107 10099 2112
<< via3 >>
rect 30308 41312 30508 41512
rect 25382 38560 25582 38760
rect 842 37854 1044 37859
rect 842 37652 847 37854
rect 847 37652 1044 37854
rect 842 37647 1044 37652
rect 30372 35654 30572 35854
rect 9051 5923 9349 5927
rect 9051 5633 9055 5923
rect 9055 5633 9345 5923
rect 9345 5633 9349 5923
rect 9051 5629 9349 5633
rect 12454 4096 12726 4100
rect 12454 3832 12458 4096
rect 12458 3832 12722 4096
rect 12722 3832 12726 4096
rect 12454 3828 12726 3832
rect 10256 3745 10519 3749
rect 10256 3490 10260 3745
rect 10260 3490 10515 3745
rect 10515 3490 10519 3745
rect 10256 3486 10519 3490
rect 9801 2407 10099 2411
rect 9801 2117 9805 2407
rect 9805 2117 10095 2407
rect 10095 2117 10099 2407
rect 9801 2113 10099 2117
<< metal4 >>
rect 798 44678 858 45152
rect 1534 44678 1594 45152
rect 2270 44678 2330 45152
rect 3006 44678 3066 45152
rect 3742 44678 3802 45152
rect 4478 44678 4538 45152
rect 5214 44678 5274 45152
rect 5950 44678 6010 45152
rect 6686 44678 6746 45152
rect 7422 44678 7482 45152
rect 8158 44678 8218 45152
rect 8894 44678 8954 45152
rect 9630 44678 9690 45152
rect 10366 44678 10426 45152
rect 11102 44678 11162 45152
rect 11838 44678 11898 45152
rect 12574 44678 12634 45152
rect 13310 44678 13370 45152
rect 14046 44678 14106 45152
rect 14782 44678 14842 45152
rect 15518 44678 15578 45152
rect 16254 44678 16314 45152
rect 16990 44678 17050 45152
rect 17726 44678 17786 45152
rect 18462 44952 18522 45152
rect 19198 44952 19258 45152
rect 19934 44952 19994 45152
rect 20670 44952 20730 45152
rect 21406 44952 21466 45152
rect 22142 44952 22202 45152
rect 22878 44952 22938 45152
rect 23614 44952 23674 45152
rect 24350 44952 24410 45152
rect 25086 44952 25146 45152
rect 25822 44952 25882 45152
rect 26558 44952 26618 45152
rect 27294 44952 27354 45152
rect 28030 44952 28090 45152
rect 28766 44952 28826 45152
rect 677 44464 17946 44678
rect 200 37854 500 44152
rect 9800 38760 10100 44152
rect 29422 41512 29622 45152
rect 30238 44952 30298 45152
rect 30974 44952 31034 45152
rect 31710 44952 31770 45152
rect 30307 41512 30509 41513
rect 29422 41312 30308 41512
rect 30508 41312 30509 41512
rect 30307 41311 30509 41312
rect 25381 38760 25583 38761
rect 9800 38560 25382 38760
rect 25582 38560 25583 38760
rect 841 37859 1045 37860
rect 841 37854 842 37859
rect 200 37652 842 37854
rect 200 7520 500 37652
rect 841 37647 842 37652
rect 1044 37647 1045 37859
rect 841 37646 1045 37647
rect 200 7220 8674 7520
rect 200 1000 500 7220
rect 8374 5928 8674 7220
rect 8374 5927 9350 5928
rect 8374 5629 9051 5927
rect 9349 5629 9350 5927
rect 8374 5628 9350 5629
rect 9800 2411 10100 38560
rect 25381 38559 25583 38560
rect 30371 35854 30573 35855
rect 30371 35654 30372 35854
rect 30572 35654 30573 35854
rect 30371 35653 30573 35654
rect 12453 4100 12727 4101
rect 12453 3828 12454 4100
rect 12726 3828 12727 4100
rect 9800 2113 9801 2411
rect 10099 2113 10100 2411
rect 9800 462 10100 2113
rect 10255 3749 10520 3750
rect 10255 3486 10256 3749
rect 10519 3486 10520 3749
rect 10255 273 10520 3486
rect 400 0 520 200
rect 4816 0 4936 200
rect 9160 120 10520 273
rect 12453 277 12727 3828
rect 30372 644 30572 35653
rect 30372 444 31412 644
rect 12453 120 13845 277
rect 31212 228 31412 444
rect 9158 0 10520 120
rect 12452 0 13846 120
rect 18064 0 18184 200
rect 22480 0 22600 200
rect 26896 0 27016 200
rect 31200 0 31432 228
use analog_mux  analog_mux_0 ~/Desktop/TinyTapeout/TinyTapeoutAnalog/tt06-programmable-thing/mag
timestamp 1713456355
transform 0 1 26232 -1 0 40002
box -240 -16 3910 4523
use inverter  inverter_0 ~/Desktop/TinyTapeout/TinyTapeoutAnalog/tt06-programmable-thing/mag
timestamp 1713454966
transform 1 0 11228 0 1 864
box -560 20 1088 6242
<< labels >>
flabel metal4 s 30974 44952 31034 45152 0 FreeSans 480 90 0 0 clk
port 0 nsew signal input
flabel metal4 s 31710 44952 31770 45152 0 FreeSans 480 90 0 0 ena
port 1 nsew signal input
flabel metal4 s 30238 44952 30298 45152 0 FreeSans 480 90 0 0 rst_n
port 2 nsew signal input
flabel metal4 s 31312 0 31432 200 0 FreeSans 960 0 0 0 ua[0]
port 3 nsew signal bidirectional
flabel metal4 s 26896 0 27016 200 0 FreeSans 960 0 0 0 ua[1]
port 4 nsew signal bidirectional
flabel metal4 s 22480 0 22600 200 0 FreeSans 960 0 0 0 ua[2]
port 5 nsew signal bidirectional
flabel metal4 s 18064 0 18184 200 0 FreeSans 960 0 0 0 ua[3]
port 6 nsew signal bidirectional
flabel metal4 s 13648 0 13768 200 0 FreeSans 960 0 0 0 ua[4]
port 7 nsew signal bidirectional
flabel metal4 s 9232 0 9352 200 0 FreeSans 960 0 0 0 ua[5]
port 8 nsew signal bidirectional
flabel metal4 s 4816 0 4936 200 0 FreeSans 960 0 0 0 ua[6]
port 9 nsew signal bidirectional
flabel metal4 s 400 0 520 200 0 FreeSans 960 0 0 0 ua[7]
port 10 nsew signal bidirectional
flabel metal4 s 29502 44952 29562 45152 0 FreeSans 480 90 0 0 ui_in[0]
port 11 nsew signal input
flabel metal4 s 28766 44952 28826 45152 0 FreeSans 480 90 0 0 ui_in[1]
port 12 nsew signal input
flabel metal4 s 28030 44952 28090 45152 0 FreeSans 480 90 0 0 ui_in[2]
port 13 nsew signal input
flabel metal4 s 27294 44952 27354 45152 0 FreeSans 480 90 0 0 ui_in[3]
port 14 nsew signal input
flabel metal4 s 26558 44952 26618 45152 0 FreeSans 480 90 0 0 ui_in[4]
port 15 nsew signal input
flabel metal4 s 25822 44952 25882 45152 0 FreeSans 480 90 0 0 ui_in[5]
port 16 nsew signal input
flabel metal4 s 25086 44952 25146 45152 0 FreeSans 480 90 0 0 ui_in[6]
port 17 nsew signal input
flabel metal4 s 24350 44952 24410 45152 0 FreeSans 480 90 0 0 ui_in[7]
port 18 nsew signal input
flabel metal4 s 23614 44952 23674 45152 0 FreeSans 480 90 0 0 uio_in[0]
port 19 nsew signal input
flabel metal4 s 22878 44952 22938 45152 0 FreeSans 480 90 0 0 uio_in[1]
port 20 nsew signal input
flabel metal4 s 22142 44952 22202 45152 0 FreeSans 480 90 0 0 uio_in[2]
port 21 nsew signal input
flabel metal4 s 21406 44952 21466 45152 0 FreeSans 480 90 0 0 uio_in[3]
port 22 nsew signal input
flabel metal4 s 20670 44952 20730 45152 0 FreeSans 480 90 0 0 uio_in[4]
port 23 nsew signal input
flabel metal4 s 19934 44952 19994 45152 0 FreeSans 480 90 0 0 uio_in[5]
port 24 nsew signal input
flabel metal4 s 19198 44952 19258 45152 0 FreeSans 480 90 0 0 uio_in[6]
port 25 nsew signal input
flabel metal4 s 18462 44952 18522 45152 0 FreeSans 480 90 0 0 uio_in[7]
port 26 nsew signal input
flabel metal4 s 5950 44952 6010 45152 0 FreeSans 480 90 0 0 uio_oe[0]
port 27 nsew signal output
flabel metal4 s 5214 44952 5274 45152 0 FreeSans 480 90 0 0 uio_oe[1]
port 28 nsew signal output
flabel metal4 s 4478 44952 4538 45152 0 FreeSans 480 90 0 0 uio_oe[2]
port 29 nsew signal output
flabel metal4 s 3742 44952 3802 45152 0 FreeSans 480 90 0 0 uio_oe[3]
port 30 nsew signal output
flabel metal4 s 3006 44952 3066 45152 0 FreeSans 480 90 0 0 uio_oe[4]
port 31 nsew signal output
flabel metal4 s 2270 44952 2330 45152 0 FreeSans 480 90 0 0 uio_oe[5]
port 32 nsew signal output
flabel metal4 s 1534 44952 1594 45152 0 FreeSans 480 90 0 0 uio_oe[6]
port 33 nsew signal output
flabel metal4 s 798 44952 858 45152 0 FreeSans 480 90 0 0 uio_oe[7]
port 34 nsew signal output
flabel metal4 s 11838 44952 11898 45152 0 FreeSans 480 90 0 0 uio_out[0]
port 35 nsew signal output
flabel metal4 s 11102 44952 11162 45152 0 FreeSans 480 90 0 0 uio_out[1]
port 36 nsew signal output
flabel metal4 s 10366 44952 10426 45152 0 FreeSans 480 90 0 0 uio_out[2]
port 37 nsew signal output
flabel metal4 s 9630 44952 9690 45152 0 FreeSans 480 90 0 0 uio_out[3]
port 38 nsew signal output
flabel metal4 s 8894 44952 8954 45152 0 FreeSans 480 90 0 0 uio_out[4]
port 39 nsew signal output
flabel metal4 s 8158 44952 8218 45152 0 FreeSans 480 90 0 0 uio_out[5]
port 40 nsew signal output
flabel metal4 s 7422 44952 7482 45152 0 FreeSans 480 90 0 0 uio_out[6]
port 41 nsew signal output
flabel metal4 s 6686 44952 6746 45152 0 FreeSans 480 90 0 0 uio_out[7]
port 42 nsew signal output
flabel metal4 s 17726 44952 17786 45152 0 FreeSans 480 90 0 0 uo_out[0]
port 43 nsew signal output
flabel metal4 s 16990 44952 17050 45152 0 FreeSans 480 90 0 0 uo_out[1]
port 44 nsew signal output
flabel metal4 s 16254 44952 16314 45152 0 FreeSans 480 90 0 0 uo_out[2]
port 45 nsew signal output
flabel metal4 s 15518 44952 15578 45152 0 FreeSans 480 90 0 0 uo_out[3]
port 46 nsew signal output
flabel metal4 s 14782 44952 14842 45152 0 FreeSans 480 90 0 0 uo_out[4]
port 47 nsew signal output
flabel metal4 s 14046 44952 14106 45152 0 FreeSans 480 90 0 0 uo_out[5]
port 48 nsew signal output
flabel metal4 s 13310 44952 13370 45152 0 FreeSans 480 90 0 0 uo_out[6]
port 49 nsew signal output
flabel metal4 s 12574 44952 12634 45152 0 FreeSans 480 90 0 0 uo_out[7]
port 50 nsew signal output
flabel metal4 200 1000 500 44152 1 FreeSans 2 0 0 0 VPWR
port 51 nsew power bidirectional
flabel metal4 9800 1000 10100 44152 1 FreeSans 2 0 0 0 VGND
port 52 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 32200 45152
<< end >>
