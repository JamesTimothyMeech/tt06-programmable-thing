magic
tech sky130A
magscale 1 2
timestamp 1713456355
<< pwell >>
rect 106 -10 382 262
<< locali >>
rect 120 4332 3560 4352
rect 120 4132 140 4332
rect 340 4156 3560 4332
rect 340 4132 400 4156
rect 120 4122 400 4132
rect 3540 4122 3560 4156
rect 120 4112 3560 4122
rect 120 4020 2420 4112
rect 1262 3942 2420 4020
rect 120 2592 944 2664
rect 120 2582 3560 2592
rect 120 2548 140 2582
rect 3280 2572 3560 2582
rect 3280 2548 3340 2572
rect 120 2396 3340 2548
rect 120 2362 140 2396
rect 3280 2372 3340 2396
rect 3540 2372 3560 2572
rect 3280 2362 3560 2372
rect 120 2268 3560 2362
<< viali >>
rect 140 4132 340 4332
rect 400 4122 3540 4156
rect 140 2548 3280 2582
rect 140 2362 3280 2396
rect 3340 2372 3540 2572
rect 100 382 134 520
<< metal1 >>
rect -166 4308 -160 4368
rect -100 4308 -94 4368
rect 120 4332 3560 4352
rect -160 4276 -100 4308
rect -240 4076 -40 4276
rect 120 4132 140 4332
rect 340 4156 598 4332
rect 650 4156 3560 4332
rect 340 4132 400 4156
rect 120 4122 400 4132
rect 3540 4122 3560 4156
rect 120 4112 3560 4122
rect 190 3912 378 3962
rect 506 3912 694 3962
rect 190 3552 236 3912
rect 282 3876 334 3882
rect 282 3582 334 3588
rect 364 3876 416 3882
rect 364 3582 416 3588
rect 506 3552 552 3912
rect 598 3876 650 3882
rect 598 3582 650 3588
rect 680 3876 732 3882
rect 680 3582 732 3588
rect 1274 3834 2256 3880
rect 190 3502 378 3552
rect 506 3502 694 3552
rect 190 3388 236 3502
rect 184 3382 242 3388
rect 506 3384 552 3502
rect 1274 3384 1320 3834
rect 1366 3796 1420 3802
rect 184 3316 242 3322
rect 502 3378 556 3384
rect 502 3320 556 3326
rect 1270 3378 1324 3384
rect 1270 3320 1324 3326
rect 190 3202 236 3316
rect 506 3202 552 3320
rect 86 3152 380 3202
rect 506 3152 800 3202
rect 86 2774 132 3152
rect 178 3108 230 3114
rect 178 2812 230 2818
rect 270 3108 324 3114
rect 270 2812 324 2818
rect 364 3108 416 3114
rect 364 2812 416 2818
rect 506 2774 552 3152
rect 598 3108 650 3114
rect 598 2812 650 2818
rect 690 3108 744 3114
rect 690 2812 744 2818
rect 784 3108 836 3114
rect 1274 2870 1320 3320
rect 1366 2902 1420 2908
rect 1494 3796 1548 3802
rect 1494 2902 1548 2908
rect 1622 3796 1676 3802
rect 1622 2902 1676 2908
rect 1750 3796 1804 3802
rect 1750 2902 1804 2908
rect 1878 3796 1932 3802
rect 1878 2902 1932 2908
rect 2006 3796 2060 3802
rect 2006 2902 2060 2908
rect 2134 3796 2188 3802
rect 2134 2902 2188 2908
rect 2262 3796 2316 3802
rect 2262 2902 2316 2908
rect 1274 2824 2256 2870
rect 3704 2842 3904 2848
rect 784 2812 836 2818
rect 86 2724 380 2774
rect 506 2724 800 2774
rect 120 2582 3560 2592
rect 120 2548 140 2582
rect 3280 2572 3560 2582
rect 3280 2548 3340 2572
rect 120 2396 178 2548
rect 230 2396 364 2548
rect 416 2396 598 2548
rect 650 2396 784 2548
rect 836 2396 3340 2548
rect 120 2362 140 2396
rect 3280 2372 3340 2396
rect 3540 2372 3560 2572
rect 3704 2556 3904 2642
rect 3280 2362 3560 2372
rect 120 2352 3560 2362
rect 3698 2442 3904 2556
rect 3698 2356 3898 2442
rect 270 2302 324 2308
rect 270 2206 324 2250
rect 270 2160 3044 2206
rect 270 1178 316 2160
rect 362 2114 416 2120
rect 362 1218 416 1232
rect 490 1978 544 2120
rect 490 1218 544 1224
rect 618 2114 672 2120
rect 618 1218 672 1360
rect 746 1978 800 2120
rect 746 1218 800 1224
rect 874 2114 928 2120
rect 874 1218 928 1360
rect 1002 1978 1056 2120
rect 1002 1218 1056 1224
rect 1130 2114 1184 2120
rect 1130 1218 1184 1360
rect 1258 1978 1312 2120
rect 1258 1218 1312 1224
rect 1386 2114 1440 2120
rect 1386 1218 1440 1360
rect 1514 1978 1568 2120
rect 1514 1218 1568 1224
rect 1642 2114 1696 2120
rect 1642 1218 1696 1360
rect 1770 1978 1824 2120
rect 1770 1218 1824 1224
rect 1898 2114 1952 2120
rect 1898 1218 1952 1360
rect 2026 1978 2080 2120
rect 2026 1218 2080 1224
rect 2154 2114 2208 2120
rect 2154 1218 2208 1360
rect 2282 1978 2336 2120
rect 2282 1218 2336 1224
rect 2410 2114 2464 2120
rect 2410 1218 2464 1360
rect 2538 1978 2592 2120
rect 2538 1218 2592 1224
rect 2666 2114 2720 2120
rect 2666 1218 2720 1360
rect 2794 1978 2848 2120
rect 2794 1218 2848 1224
rect 2922 2114 2976 2120
rect 2922 1218 2976 1360
rect 3050 2114 3104 2120
rect 3050 1218 3104 1224
rect 270 1132 3044 1178
rect 2666 972 3098 996
rect 2666 912 2696 972
rect 3068 912 3098 972
rect 54 520 798 646
rect 54 382 100 520
rect 134 382 798 520
rect 2666 414 3098 912
rect 54 252 798 382
rect 54 244 120 252
rect 106 12 120 244
rect 360 244 798 252
rect 360 184 382 244
rect 360 12 1442 184
rect 106 -16 1442 12
rect 2148 0 2473 202
rect 2675 0 2681 202
<< via1 >>
rect -160 4308 -100 4368
rect 140 4132 340 4332
rect 598 4156 650 4332
rect 598 4132 650 4156
rect 282 3588 334 3876
rect 364 3588 416 3876
rect 598 3588 650 3876
rect 680 3588 732 3876
rect 184 3322 242 3382
rect 502 3326 556 3378
rect 1270 3326 1324 3378
rect 178 2818 230 3108
rect 270 2818 324 3108
rect 364 2818 416 3108
rect 598 2818 650 3108
rect 690 2818 744 3108
rect 784 2818 836 3108
rect 1366 2908 1420 3796
rect 1494 2908 1548 3796
rect 1622 2908 1676 3796
rect 1750 2908 1804 3796
rect 1878 2908 1932 3796
rect 2006 2908 2060 3796
rect 2134 2908 2188 3796
rect 2262 2908 2316 3796
rect 3704 2642 3904 2842
rect 178 2548 230 2572
rect 364 2548 416 2572
rect 598 2548 650 2572
rect 784 2548 836 2572
rect 178 2396 230 2548
rect 364 2396 416 2548
rect 598 2396 650 2548
rect 784 2396 836 2548
rect 178 2372 230 2396
rect 364 2372 416 2396
rect 598 2372 650 2396
rect 784 2372 836 2396
rect 3340 2372 3540 2572
rect 270 2250 324 2302
rect 362 1232 416 2114
rect 490 1224 544 1978
rect 618 1360 672 2114
rect 746 1224 800 1978
rect 874 1360 928 2114
rect 1002 1224 1056 1978
rect 1130 1360 1184 2114
rect 1258 1224 1312 1978
rect 1386 1360 1440 2114
rect 1514 1224 1568 1978
rect 1642 1360 1696 2114
rect 1770 1224 1824 1978
rect 1898 1360 1952 2114
rect 2026 1224 2080 1978
rect 2154 1360 2208 2114
rect 2282 1224 2336 1978
rect 2410 1360 2464 2114
rect 2538 1224 2592 1978
rect 2666 1360 2720 2114
rect 2794 1224 2848 1978
rect 2922 1360 2976 2114
rect 3050 1224 3104 2114
rect 2696 912 3068 972
rect 120 12 360 252
rect 2473 0 2675 202
<< metal2 >>
rect -160 4518 -100 4520
rect -167 4462 -158 4518
rect -102 4462 -93 4518
rect -160 4368 -100 4462
rect -160 4302 -100 4308
rect 120 4332 360 4352
rect 120 4132 140 4332
rect 340 4132 360 4332
rect 120 4112 360 4132
rect 598 4332 650 4352
rect 282 3876 334 4112
rect 282 3582 334 3588
rect 364 3876 416 3882
rect 184 3382 242 3392
rect 364 3372 416 3588
rect 598 3876 650 4132
rect 1650 4342 2050 4352
rect 1650 4062 1756 4342
rect 1366 3962 1756 4062
rect 1924 4062 2050 4342
rect 1924 4026 2190 4062
rect 1924 3962 2188 4026
rect 598 3582 650 3588
rect 680 3876 732 3882
rect 496 3372 502 3378
rect 184 3312 242 3322
rect 270 3332 502 3372
rect 178 3108 230 3114
rect 178 2572 230 2818
rect 178 2352 230 2372
rect 270 3108 324 3332
rect 496 3326 502 3332
rect 556 3326 562 3378
rect 680 3372 732 3588
rect 1366 3862 2188 3962
rect 1366 3796 1420 3862
rect 1264 3372 1270 3378
rect 680 3332 1270 3372
rect 270 2302 324 2818
rect 364 3108 416 3114
rect 364 2572 416 2818
rect 364 2352 416 2372
rect 598 3108 650 3114
rect 598 2572 650 2818
rect 690 3108 744 3332
rect 1264 3326 1270 3332
rect 1324 3326 1330 3378
rect 690 2812 744 2818
rect 784 3108 836 3114
rect 1366 2902 1420 2908
rect 1494 3796 1548 3802
rect 598 2352 650 2372
rect 784 2572 836 2818
rect 1494 2842 1548 2908
rect 1622 3796 1676 3862
rect 1622 2902 1676 2908
rect 1750 3796 1804 3802
rect 1750 2842 1804 2908
rect 1878 3796 1932 3862
rect 1878 2902 1932 2908
rect 2006 3796 2060 3802
rect 2006 2842 2060 2908
rect 2134 3796 2188 3862
rect 2134 2902 2188 2908
rect 2262 3796 2316 3802
rect 2262 2842 2316 2908
rect 1494 2742 3704 2842
rect 1494 2642 1756 2742
rect 784 2352 836 2372
rect 1640 2362 1756 2642
rect 1924 2642 3704 2742
rect 3904 2642 3910 2842
rect 1924 2362 2040 2642
rect 1640 2252 2040 2362
rect 3320 2572 3560 2592
rect 3320 2372 3340 2572
rect 3540 2372 3560 2572
rect 3320 2352 3560 2372
rect 270 2244 324 2250
rect 416 2120 2922 2252
rect 3050 2166 3450 2176
rect 362 2114 2978 2120
rect 416 2052 618 2114
rect 362 1218 416 1232
rect 490 1978 544 1984
rect 672 2052 874 2114
rect 618 1354 672 1360
rect 746 1978 800 1984
rect 544 1224 746 1286
rect 928 2052 1130 2114
rect 874 1354 928 1360
rect 1002 1978 1056 1984
rect 800 1224 1002 1286
rect 1184 2052 1386 2114
rect 1130 1354 1184 1360
rect 1258 1978 1312 1984
rect 1056 1224 1258 1286
rect 1440 2052 1642 2114
rect 1386 1354 1440 1360
rect 1514 1978 1568 1984
rect 1312 1224 1514 1286
rect 1696 2052 1898 2114
rect 1642 1354 1696 1360
rect 1770 1978 1824 1984
rect 1568 1224 1770 1286
rect 1952 2052 2154 2114
rect 1898 1354 1952 1360
rect 2026 1978 2080 1984
rect 1824 1224 2026 1286
rect 2208 2052 2410 2114
rect 2154 1354 2208 1360
rect 2282 1978 2336 1984
rect 2080 1224 2282 1286
rect 2464 2052 2666 2114
rect 2410 1354 2464 1360
rect 2538 1978 2592 1984
rect 2336 1224 2538 1286
rect 2720 2052 2922 2114
rect 2666 1354 2720 1360
rect 2794 1978 2848 1984
rect 2592 1224 2794 1286
rect 2976 2052 2978 2114
rect 3050 2114 3056 2166
rect 2922 1354 2976 1360
rect 3344 1914 3450 2166
rect 2848 1224 3050 1286
rect 3104 1224 3450 1914
rect 490 1086 3450 1224
rect 1458 972 3450 1086
rect 1458 912 2696 972
rect 3068 912 3450 972
rect 1458 886 3450 912
rect 125 252 355 256
rect 114 12 120 252
rect 360 12 366 252
rect 2473 202 2675 208
rect 125 8 355 12
rect 2675 0 2719 202
rect 2921 0 2930 202
rect 2473 -6 2675 0
<< via2 >>
rect -158 4462 -102 4518
rect 140 4132 340 4332
rect 184 3322 242 3382
rect 1756 3962 1924 4342
rect 1756 2362 1924 2742
rect 3340 2372 3540 2572
rect 3056 2114 3344 2166
rect 3056 1914 3104 2114
rect 3104 1914 3344 2114
rect 125 17 355 247
rect 2719 0 2921 202
<< metal3 >>
rect -163 4520 -97 4523
rect -163 4518 950 4520
rect -163 4462 -158 4518
rect -102 4462 950 4518
rect -163 4460 950 4462
rect -163 4457 -97 4460
rect 120 4332 360 4352
rect 120 4132 140 4332
rect 340 4132 360 4332
rect 120 4112 360 4132
rect 178 3382 248 3388
rect 890 3382 950 4460
rect 1750 4346 1930 4352
rect 1750 3958 1756 4346
rect 1924 4132 1930 4346
rect 1924 3958 3140 4132
rect 1750 3952 3140 3958
rect 178 3322 184 3382
rect 242 3322 950 3382
rect 178 3316 248 3322
rect 1750 2746 1930 2752
rect 1750 2358 1756 2746
rect 1924 2358 1930 2746
rect 1750 2352 1930 2358
rect 2960 2172 3140 3952
rect 3320 2572 3560 2592
rect 3320 2372 3340 2572
rect 3540 2372 3560 2572
rect 3320 2352 3560 2372
rect 2960 2166 3350 2172
rect 2960 1914 3056 2166
rect 3344 1914 3350 2166
rect 2960 1908 3350 1914
rect 121 252 359 257
rect 120 251 360 252
rect 120 13 121 251
rect 359 13 360 251
rect 120 12 360 13
rect 2714 202 2926 207
rect 121 7 359 12
rect 2714 0 2719 202
rect 2921 0 2965 202
rect 3167 0 3173 202
rect 2714 -5 2926 0
<< via3 >>
rect 140 4132 340 4332
rect 1756 4342 1924 4346
rect 1756 3962 1924 4342
rect 1756 3958 1924 3962
rect 1756 2742 1924 2746
rect 1756 2362 1924 2742
rect 1756 2358 1924 2362
rect 3340 2372 3540 2572
rect 121 247 359 251
rect 121 17 125 247
rect 125 17 355 247
rect 355 17 359 247
rect 121 13 359 17
rect 2965 0 3167 202
<< metal4 >>
rect 120 4332 360 4352
rect 120 4132 140 4332
rect 340 4132 360 4332
rect 120 251 360 4132
rect 1750 4346 1930 4352
rect 1750 3958 1756 4346
rect 1924 3958 1930 4346
rect 1750 3952 1930 3958
rect 1750 2746 1930 2752
rect 1750 2358 1756 2746
rect 1924 2358 1930 2746
rect 1750 2352 1930 2358
rect 3320 2572 3560 4352
rect 3320 2372 3340 2572
rect 3540 2372 3560 2572
rect 120 13 121 251
rect 359 13 360 251
rect 120 0 360 13
rect 2964 202 3168 203
rect 3320 202 3560 2372
rect 2964 0 2965 202
rect 3167 0 3560 202
rect 2964 -1 3168 0
use sky130_fd_pr__nfet_01v8_lvt_9LK66Y  sky130_fd_pr__nfet_01v8_lvt_9LK66Y_0
timestamp 1712480545
transform 1 0 1841 0 1 3352
box -615 -660 615 660
use sky130_fd_pr__nfet_01v8_NRQ53D  sky130_fd_pr__nfet_01v8_NRQ53D_0
timestamp 1712308627
transform 1 0 665 0 1 3732
box -211 -360 211 360
use sky130_fd_pr__nfet_01v8_NRQ53D  sky130_fd_pr__nfet_01v8_NRQ53D_1
timestamp 1712308627
transform 1 0 349 0 1 3732
box -211 -360 211 360
use sky130_fd_pr__pfet_01v8_lvt_MUCXQQ  sky130_fd_pr__pfet_01v8_lvt_MUCXQQ_0
timestamp 1713454966
transform 1 0 1733 0 1 1669
box -1511 -669 1511 669
use sky130_fd_pr__pfet_01v8_XJBLHL  sky130_fd_pr__pfet_01v8_XJBLHL_0
timestamp 1713454966
transform 1 0 297 0 1 2963
box -263 -369 263 369
use sky130_fd_pr__pfet_01v8_XJBLHL  sky130_fd_pr__pfet_01v8_XJBLHL_1
timestamp 1713454966
transform 1 0 717 0 1 2963
box -263 -369 263 369
use sky130_fd_pr__res_xhigh_po_0p35_KNBXRF  XR1
timestamp 1713452737
transform 0 1 1664 -1 0 451
box -201 -1598 201 1598
<< labels >>
rlabel metal4 120 0 360 4352 1 VGND
port 1 n ground input
rlabel metal4 3320 0 3560 4352 1 VPWR
port 2 n power input
rlabel metal4 1750 3952 1930 4352 1 mod
port 3 n analog bidirectional
rlabel metal4 1750 2352 1930 2752 1 bus
port 4 n analog bidirectional
rlabel metal3 890 4172 950 4352 1 ctrl
port 5 n signal input
flabel metal1 1242 -16 1442 184 0 FreeSans 256 0 0 0 VGND
flabel metal1 2150 2 2350 202 0 FreeSans 256 0 0 0 VPWR
port 0 nsew
flabel metal1 2786 674 2986 874 0 FreeSans 256 0 0 0 mod
flabel metal1 3698 2356 3898 2556 0 FreeSans 256 0 0 0 bus
flabel metal1 -240 4076 -40 4276 0 FreeSans 256 0 0 0 ctrl
<< properties >>
string FIXED_BBOX 0 0 3680 4352
<< end >>
