magic
tech sky130A
magscale 1 2
timestamp 1713204041
<< pwell >>
rect 422 448 456 2346
rect 680 432 876 2392
<< viali >>
rect 320 3940 354 5798
rect 308 462 342 2346
<< metal1 >>
rect -559 6042 678 6242
rect -559 5980 -359 6042
rect -559 5946 -358 5980
rect -559 3852 -359 5946
rect 478 5932 678 6042
rect -182 5868 214 5890
rect -182 5798 448 5868
rect -182 3940 320 5798
rect 354 3940 466 5798
rect -182 3910 256 3940
rect 314 3932 366 3940
rect 314 3930 358 3932
rect 690 3910 1088 5888
rect -559 3818 -358 3852
rect -559 3204 -359 3818
rect 480 3218 680 3858
rect -560 3202 -359 3204
rect 478 3202 682 3218
rect 890 3204 1088 3910
rect -560 3004 682 3202
rect 888 3004 1088 3204
rect -559 3002 682 3004
rect -559 220 -359 3002
rect 478 2444 682 3002
rect 890 2815 1088 3004
rect 894 2392 1087 2815
rect -182 2346 228 2392
rect 296 2346 348 2358
rect -182 462 308 2346
rect 342 462 456 2346
rect -182 448 456 462
rect -182 432 240 448
rect 680 432 1087 2392
rect -182 428 232 432
rect 468 220 668 380
rect -559 20 668 220
use sky130_fd_pr__pfet_01v8_GGAEPD  XM1
timestamp 1713203168
transform 1 0 578 0 1 4899
box -296 -1219 296 1219
use sky130_fd_pr__nfet_01v8_6WXQK8  XM2
timestamp 1713203168
transform -1 0 568 0 1 1412
box -296 -1210 296 1210
<< labels >>
flabel metal1 888 3004 1088 3204 0 FreeSans 256 0 0 0 OUT
port 2 nsew
flabel metal1 -560 3004 -360 3204 0 FreeSans 256 0 0 0 IN
port 3 nsew
flabel metal1 -176 5680 24 5880 0 FreeSans 256 0 0 0 VDD
port 0 nsew
flabel metal1 -170 440 30 640 0 FreeSans 256 0 0 0 VSS
port 1 nsew
<< end >>
