magic
tech sky130A
magscale 1 2
timestamp 1713118345
<< pwell >>
rect 422 432 456 2392
rect 680 432 876 2392
<< viali >>
rect 414 6048 742 6082
rect 320 3934 354 5856
rect 308 462 342 2362
rect 404 238 732 272
<< metal1 >>
rect -334 6216 -298 6218
rect -562 6018 -298 6216
rect 142 6082 874 6218
rect 142 6048 414 6082
rect 742 6048 874 6082
rect 142 6018 874 6048
rect -562 6016 242 6018
rect -559 5946 662 5980
rect -559 3852 -478 5946
rect -418 5878 466 5888
rect -418 4014 -306 5878
rect 151 5856 466 5878
rect 151 4014 320 5856
rect -418 3934 320 4014
rect 354 3934 466 5856
rect -418 3910 466 3934
rect 690 3910 1088 5888
rect -559 3818 662 3852
rect -559 3204 -359 3818
rect 890 3204 1088 3910
rect -560 3004 -359 3204
rect 888 3004 1088 3204
rect -559 2484 -359 3004
rect 890 2815 1088 3004
rect -559 2450 668 2484
rect -559 374 -478 2450
rect 894 2392 1087 2815
rect -422 2362 456 2392
rect -422 2289 308 2362
rect -422 432 -303 2289
rect -309 427 -303 432
rect 176 462 308 2289
rect 342 462 456 2362
rect 176 432 456 462
rect 680 432 1087 2392
rect 176 427 182 432
rect -303 419 176 427
rect -559 339 496 374
rect -559 338 -478 339
rect -308 300 -191 306
rect -91 300 178 306
rect -558 96 -308 296
rect 178 296 184 300
rect 178 272 864 296
rect 178 238 404 272
rect 732 238 864 272
rect 178 211 864 238
rect -314 94 -308 96
rect 180 96 864 211
rect 180 94 186 96
rect 732 94 864 96
rect -218 88 -212 94
rect 100 88 180 94
rect -97 86 100 88
<< via1 >>
rect -298 6018 142 6218
rect -306 4014 151 5878
rect -303 427 176 2289
rect -308 211 178 300
rect -308 94 180 211
rect -212 88 100 94
<< metal2 >>
rect -306 6218 151 6220
rect -306 6018 -298 6218
rect 142 6018 151 6218
rect -306 5878 151 6018
rect -306 4008 151 4014
rect -303 2289 176 2297
rect -309 427 -303 1363
rect 176 427 182 1363
rect -308 300 178 427
rect -314 183 -308 300
rect 178 211 184 300
rect 180 94 186 211
rect -308 88 -212 94
rect 100 88 180 94
rect -212 86 -95 88
use sky130_fd_pr__pfet_01v8_GGAEPD  XM1
timestamp 1713027578
transform 1 0 578 0 1 4899
box -296 -1219 296 1219
use sky130_fd_pr__nfet_01v8_6WXQK8  XM2
timestamp 1713027578
transform -1 0 568 0 1 1412
box -296 -1210 296 1210
<< labels >>
flabel metal1 -562 6016 -362 6216 0 FreeSans 256 0 0 0 VDD
port 0 nsew
flabel metal1 -558 96 -358 296 0 FreeSans 256 0 0 0 VSS
port 1 nsew
flabel metal1 888 3004 1088 3204 0 FreeSans 256 0 0 0 OUT
port 2 nsew
flabel metal1 -560 3004 -360 3204 0 FreeSans 256 0 0 0 IN
port 3 nsew
<< end >>
