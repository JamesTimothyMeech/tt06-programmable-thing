magic
tech sky130A
magscale 1 2
timestamp 1713480354
<< metal1 >>
rect 27952 41286 28152 41292
rect 27212 41260 27412 41266
rect 24830 41060 27212 41260
rect 24830 40906 25030 41060
rect 27212 41054 27412 41060
rect 27952 40914 28152 41086
rect 20564 40706 25030 40906
rect 25200 40714 28152 40914
rect 20564 40542 20764 40706
rect 25200 40542 25400 40714
rect 15984 40342 20764 40542
rect 20932 40342 25400 40542
rect 30308 40674 30508 40680
rect 15984 40062 16184 40342
rect 20932 40046 21132 40342
rect 25582 40240 28688 40440
rect 28888 40240 28894 40440
rect 25582 40044 25782 40240
rect 30308 40042 30508 40474
rect 12092 38960 12098 39160
rect 16816 38820 16986 39020
rect 9324 38760 9524 38766
rect 9524 38560 12072 38760
rect 21444 38560 21668 38760
rect 26126 38560 26416 38760
rect 9324 38554 9524 38560
rect 10023 37854 12110 37874
rect 1365 37652 1371 37854
rect 1573 37672 12110 37854
rect 1573 37652 10158 37672
rect 11898 37652 12045 37672
rect 16816 37652 17041 37854
rect 21444 37652 21669 37854
rect 26126 37652 26434 37854
rect 14350 36308 20184 36318
rect 14350 36304 24768 36308
rect 14350 36118 30372 36304
rect 19212 36108 30372 36118
rect 23884 36104 30372 36108
rect 30572 36104 30578 36304
rect 9392 33406 9398 33606
rect 9598 33406 12022 33606
rect 1635 32489 1641 32691
rect 1843 32489 12087 32691
rect 14242 31082 19076 31106
rect 23544 31082 28276 31122
rect 14242 30922 28276 31082
rect 14242 30906 23650 30922
rect 18964 30882 23650 30906
rect 11428 28262 11434 28462
rect 11634 28262 25956 28462
rect 1647 27354 1653 27556
rect 1855 27354 25974 27556
rect 11096 5928 11396 6474
rect 11096 5622 11396 5628
rect 12079 4101 12353 4107
rect 10249 3833 10255 4098
rect 10520 3833 10870 4098
rect 12079 3821 12353 3827
rect 11122 2412 11422 2418
rect 11122 1730 11422 2112
<< via1 >>
rect 27212 41060 27412 41260
rect 27952 41086 28152 41286
rect 30308 40474 30508 40674
rect 28688 40240 28888 40440
rect 11898 38960 12092 39160
rect 9324 38560 9524 38760
rect 1371 37652 1573 37854
rect 30372 36104 30572 36304
rect 9398 33406 9598 33606
rect 1641 32489 1843 32691
rect 11434 28262 11634 28462
rect 1653 27354 1855 27556
rect 11096 5628 11396 5928
rect 10255 3833 10520 4098
rect 12079 3827 12353 4101
rect 11122 2112 11422 2412
<< metal2 >>
rect 27952 41616 28152 41625
rect 27212 41548 27412 41557
rect 27212 41260 27412 41348
rect 27952 41286 28152 41416
rect 27206 41060 27212 41260
rect 27412 41060 27418 41260
rect 27946 41086 27952 41286
rect 28152 41086 28158 41286
rect 30308 41052 30508 41061
rect 28688 41012 28888 41021
rect 28688 40440 28888 40812
rect 30308 40674 30508 40852
rect 30302 40474 30308 40674
rect 30508 40474 30514 40674
rect 28688 40234 28888 40240
rect 11898 39160 12092 39166
rect 9324 39042 9524 39051
rect 11898 38954 12092 38960
rect 9324 38760 9524 38842
rect 9318 38560 9324 38760
rect 9524 38560 9530 38760
rect 847 37854 1049 37863
rect 1371 37854 1573 37860
rect 1049 37652 1371 37854
rect 847 37643 1049 37652
rect 1371 37646 1573 37652
rect 30372 36304 30572 36310
rect 30372 36086 30572 36104
rect 30372 35877 30572 35886
rect 25555 34792 25564 34848
rect 25620 34792 25629 34848
rect 9398 33878 9598 33887
rect 9398 33606 9598 33678
rect 9398 33400 9598 33406
rect 1641 32691 1843 32697
rect 1340 32489 1349 32691
rect 1551 32489 1641 32691
rect 1641 32483 1843 32489
rect 28364 31132 28564 31344
rect 28355 30932 28364 31132
rect 28564 30932 28573 31132
rect 11434 28462 11634 28468
rect 11425 28262 11434 28462
rect 11634 28262 11643 28462
rect 11434 28256 11634 28262
rect 1653 27556 1855 27562
rect 1644 27354 1653 27556
rect 1855 27354 1864 27556
rect 1653 27348 1855 27354
rect 28414 25994 28614 26200
rect 28405 25794 28414 25994
rect 28614 25794 28623 25994
rect 9050 5923 11096 5928
rect 9046 5633 9055 5923
rect 9345 5633 11096 5923
rect 9050 5628 11096 5633
rect 11396 5628 11402 5928
rect 10255 4098 10520 4104
rect 12458 4101 12722 4105
rect 10255 3745 10520 3833
rect 12073 3827 12079 4101
rect 12353 4096 12727 4101
rect 12353 3832 12458 4096
rect 12722 3832 12727 4096
rect 12353 3827 12727 3832
rect 12458 3823 12722 3827
rect 10251 3490 10260 3745
rect 10515 3490 10524 3745
rect 10255 3485 10520 3490
rect 9805 2412 10095 2416
rect 9800 2407 11122 2412
rect 9800 2117 9805 2407
rect 10095 2117 11122 2407
rect 9800 2112 11122 2117
rect 11422 2112 11428 2412
rect 9805 2108 10095 2112
<< via2 >>
rect 27212 41348 27412 41548
rect 27952 41416 28152 41616
rect 28688 40812 28888 41012
rect 30308 40852 30508 41052
rect 9324 38842 9524 39042
rect 847 37652 1049 37854
rect 30372 35886 30572 36086
rect 25564 34792 25620 34848
rect 9398 33678 9598 33878
rect 1349 32489 1551 32691
rect 28364 30932 28564 31132
rect 11434 28262 11634 28462
rect 1653 27354 1855 27556
rect 28414 25794 28614 25994
rect 9055 5633 9345 5923
rect 12458 3832 12722 4096
rect 10260 3490 10515 3745
rect 9805 2117 10095 2407
<< metal3 >>
rect 27952 41988 28152 41994
rect 27952 41621 28152 41788
rect 27947 41616 28157 41621
rect 27207 41553 27417 41559
rect 27947 41416 27952 41616
rect 28152 41416 28157 41616
rect 27947 41411 28157 41416
rect 30308 41512 30508 41518
rect 27207 41348 27212 41353
rect 27412 41348 27417 41353
rect 27207 41343 27417 41348
rect 28688 41314 28888 41320
rect 28688 41017 28888 41114
rect 30308 41057 30508 41312
rect 30303 41052 30513 41057
rect 28683 41012 28893 41017
rect 28683 40812 28688 41012
rect 28888 40812 28893 41012
rect 30303 40852 30308 41052
rect 30508 40852 30513 41052
rect 30303 40847 30513 40852
rect 28683 40807 28893 40812
rect 9324 39280 9524 39286
rect 9324 39047 9524 39080
rect 9319 39042 9529 39047
rect 9319 38842 9324 39042
rect 9524 38842 9529 39042
rect 9319 38837 9529 38842
rect 836 37647 842 37859
rect 1044 37854 1054 37859
rect 1049 37652 1054 37854
rect 1044 37647 1054 37652
rect 30367 36086 30577 36091
rect 30367 35886 30372 36086
rect 30572 35886 30577 36086
rect 25554 35818 25560 35882
rect 25624 35818 25630 35882
rect 30367 35881 30577 35886
rect 30372 35854 30572 35881
rect 16344 35436 16408 35442
rect 16344 35366 16408 35372
rect 16346 34626 16406 35366
rect 20980 35326 21044 35332
rect 20980 35256 21044 35262
rect 20982 34730 21042 35256
rect 25562 34853 25622 35818
rect 30174 35648 30180 35712
rect 30244 35648 30250 35712
rect 30372 35648 30572 35654
rect 25559 34848 25625 34853
rect 30182 34850 30242 35648
rect 25559 34792 25564 34848
rect 25620 34792 25625 34848
rect 25559 34787 25625 34792
rect 25562 34620 25622 34787
rect 9393 33883 9603 33889
rect 9393 33678 9398 33683
rect 9598 33678 9603 33683
rect 9393 33673 9603 33678
rect 1344 32691 1556 32696
rect 995 32489 1001 32691
rect 1203 32489 1349 32691
rect 1551 32489 1556 32691
rect 1344 32484 1556 32489
rect 28359 31132 28569 31137
rect 28359 30932 28364 31132
rect 28564 30932 29782 31132
rect 29982 30932 29988 31132
rect 28359 30927 28569 30932
rect 30230 30360 30294 30366
rect 30230 30290 30294 30296
rect 30232 29592 30292 30290
rect 11423 28257 11429 28467
rect 11629 28462 11639 28467
rect 11634 28262 11639 28462
rect 11629 28257 11639 28262
rect 1648 27556 1860 27561
rect 1163 27354 1169 27556
rect 1371 27354 1653 27556
rect 1855 27354 1860 27556
rect 1648 27349 1860 27354
rect 28409 25994 28619 25999
rect 29432 25994 29632 26000
rect 28409 25794 28414 25994
rect 28614 25794 29432 25994
rect 28409 25789 28619 25794
rect 29432 25788 29632 25794
rect 9051 5928 9349 5933
rect 9050 5927 9350 5928
rect 9050 5629 9051 5927
rect 9349 5629 9350 5927
rect 9050 5628 9350 5629
rect 9051 5623 9349 5628
rect 12453 4100 12727 4101
rect 12448 3828 12454 4100
rect 12726 3828 12732 4100
rect 12453 3827 12727 3828
rect 10255 3749 10520 3750
rect 10250 3486 10256 3749
rect 10519 3486 10525 3749
rect 10255 3485 10520 3486
rect 9801 2412 10099 2417
rect 9800 2411 10100 2412
rect 9800 2113 9801 2411
rect 10099 2113 10100 2411
rect 9800 2112 10100 2113
rect 9801 2107 10099 2112
<< via3 >>
rect 27952 41788 28152 41988
rect 27207 41548 27417 41553
rect 27207 41353 27212 41548
rect 27212 41353 27412 41548
rect 27412 41353 27417 41548
rect 28688 41114 28888 41314
rect 30308 41312 30508 41512
rect 9324 39080 9524 39280
rect 842 37854 1044 37859
rect 842 37652 847 37854
rect 847 37652 1044 37854
rect 842 37647 1044 37652
rect 25560 35818 25624 35882
rect 16344 35372 16408 35436
rect 20980 35262 21044 35326
rect 30180 35648 30244 35712
rect 30372 35654 30572 35854
rect 9393 33878 9603 33883
rect 9393 33683 9398 33878
rect 9398 33683 9598 33878
rect 9598 33683 9603 33878
rect 1001 32489 1203 32691
rect 29782 30932 29982 31132
rect 30230 30296 30294 30360
rect 11429 28462 11629 28467
rect 11429 28262 11434 28462
rect 11434 28262 11629 28462
rect 11429 28257 11629 28262
rect 1169 27354 1371 27556
rect 29432 25794 29632 25994
rect 9051 5923 9349 5927
rect 9051 5633 9055 5923
rect 9055 5633 9345 5923
rect 9345 5633 9349 5923
rect 9051 5629 9349 5633
rect 12454 4096 12726 4100
rect 12454 3832 12458 4096
rect 12458 3832 12722 4096
rect 12722 3832 12726 4096
rect 12454 3828 12726 3832
rect 10256 3745 10519 3749
rect 10256 3490 10260 3745
rect 10260 3490 10515 3745
rect 10515 3490 10519 3745
rect 10256 3486 10519 3490
rect 9801 2407 10099 2411
rect 9801 2117 9805 2407
rect 9805 2117 10095 2407
rect 10095 2117 10099 2407
rect 9801 2113 10099 2117
<< metal4 >>
rect 798 44678 858 45152
rect 1534 44678 1594 45152
rect 2270 44678 2330 45152
rect 3006 44678 3066 45152
rect 3742 44678 3802 45152
rect 4478 44678 4538 45152
rect 5214 44678 5274 45152
rect 5950 44678 6010 45152
rect 6686 44678 6746 45152
rect 7422 44678 7482 45152
rect 8158 44678 8218 45152
rect 8894 44678 8954 45152
rect 9630 44678 9690 45152
rect 10366 44678 10426 45152
rect 11102 44678 11162 45152
rect 11838 44678 11898 45152
rect 12574 44678 12634 45152
rect 13310 44678 13370 45152
rect 14046 44678 14106 45152
rect 14782 44678 14842 45152
rect 15518 44678 15578 45152
rect 16254 44678 16314 45152
rect 16990 44678 17050 45152
rect 17726 44678 17786 45152
rect 18462 44952 18522 45152
rect 19198 44952 19258 45152
rect 19934 44952 19994 45152
rect 20670 44952 20730 45152
rect 21406 44952 21466 45152
rect 22142 44952 22202 45152
rect 22878 44952 22938 45152
rect 677 44464 17946 44678
rect 11834 44460 11898 44464
rect 200 37854 500 44152
rect 9323 39280 9525 39281
rect 9800 39280 10100 44152
rect 23614 41636 23674 45152
rect 24350 41832 24410 45152
rect 19886 41576 23674 41636
rect 24276 41772 24410 41832
rect 9323 39080 9324 39280
rect 9524 39080 10100 39280
rect 9323 39079 9525 39080
rect 9800 38760 10100 39080
rect 9800 38560 10158 38760
rect 841 37859 1045 37860
rect 841 37854 842 37859
rect 200 37652 842 37854
rect 200 32691 500 37652
rect 841 37647 842 37652
rect 1044 37647 1045 37859
rect 841 37646 1045 37647
rect 9392 33883 9604 33884
rect 9800 33883 10100 38560
rect 9392 33683 9393 33883
rect 9603 33683 10100 33883
rect 9392 33682 9604 33683
rect 9800 33606 10100 33683
rect 9800 33406 10104 33606
rect 1000 32691 1204 32692
rect 200 32489 1001 32691
rect 1203 32489 1204 32691
rect 200 27556 500 32489
rect 1000 32488 1204 32489
rect 9800 28462 10100 33406
rect 10580 30192 10640 41374
rect 10802 30382 10862 41374
rect 11102 40830 11162 41374
rect 19886 41286 19946 41576
rect 24276 41496 24336 41772
rect 25086 41696 25146 45152
rect 11016 40770 11162 40830
rect 15302 41226 19946 41286
rect 20030 41436 24336 41496
rect 24436 41636 25146 41696
rect 11016 30568 11076 40770
rect 11834 40688 11898 40690
rect 11186 40672 11898 40688
rect 15302 40672 15362 41226
rect 20030 41150 20090 41436
rect 24436 41354 24496 41636
rect 25822 41536 25882 45152
rect 11186 40624 15362 40672
rect 11186 30742 11250 40624
rect 11844 40612 15362 40624
rect 15436 41090 20090 41150
rect 20172 41294 24496 41354
rect 24570 41476 25882 41536
rect 15436 40542 15496 41090
rect 20172 41010 20232 41294
rect 24570 41198 24630 41476
rect 26558 41394 26618 45152
rect 27212 41554 27412 45152
rect 27951 45030 28152 45152
rect 27952 41989 28152 45030
rect 27951 41988 28153 41989
rect 27951 41788 27952 41988
rect 28152 41788 28153 41988
rect 27951 41787 28153 41788
rect 11322 40482 15496 40542
rect 15566 40950 20232 41010
rect 20304 41138 24630 41198
rect 24712 41334 26618 41394
rect 27206 41553 27418 41554
rect 27206 41353 27207 41553
rect 27417 41353 27418 41553
rect 27206 41352 27418 41353
rect 11322 35614 11382 40482
rect 15566 40406 15626 40950
rect 20304 40854 20364 41138
rect 24712 41074 24772 41334
rect 28688 41315 28888 45152
rect 29422 41512 29622 45152
rect 30238 44952 30298 45152
rect 30974 44952 31034 45152
rect 31710 44952 31770 45152
rect 30307 41512 30509 41513
rect 28687 41314 28889 41315
rect 28687 41114 28688 41314
rect 28888 41114 28889 41314
rect 29422 41312 30308 41512
rect 30508 41312 30509 41512
rect 30307 41311 30509 41312
rect 28687 41113 28889 41114
rect 11454 40346 15626 40406
rect 15728 40794 20364 40854
rect 20432 41014 24772 41074
rect 11454 35734 11514 40346
rect 15728 40246 15788 40794
rect 20432 40700 20492 41014
rect 11584 40186 15788 40246
rect 15860 40640 20492 40700
rect 11584 35882 11644 40186
rect 15860 40098 15920 40640
rect 11726 40038 15920 40098
rect 11726 36006 11786 40038
rect 16030 39646 17840 39886
rect 20944 39644 22520 39884
rect 25022 39644 26498 39884
rect 15226 36446 17436 36686
rect 20214 36444 22064 36684
rect 25356 36444 26680 36684
rect 11726 35946 30242 36006
rect 25559 35882 25625 35883
rect 11584 35880 25206 35882
rect 25559 35880 25560 35882
rect 11584 35822 25560 35880
rect 25136 35820 25560 35822
rect 25559 35818 25560 35820
rect 25624 35818 25625 35882
rect 25559 35817 25625 35818
rect 11454 35674 21042 35734
rect 30182 35713 30242 35946
rect 30371 35854 30573 35855
rect 11322 35612 16096 35614
rect 11322 35554 16406 35612
rect 16046 35552 16406 35554
rect 16346 35437 16406 35552
rect 16343 35436 16409 35437
rect 16343 35372 16344 35436
rect 16408 35372 16409 35436
rect 16343 35371 16409 35372
rect 20982 35327 21042 35674
rect 30179 35712 30245 35713
rect 30179 35648 30180 35712
rect 30244 35648 30245 35712
rect 30371 35654 30372 35854
rect 30572 35654 30573 35854
rect 30371 35653 30573 35654
rect 30179 35647 30245 35648
rect 20979 35326 21045 35327
rect 20979 35262 20980 35326
rect 21044 35262 21045 35326
rect 20979 35261 21045 35262
rect 16008 34426 17530 34666
rect 20646 34466 22024 34706
rect 25232 34488 26716 34728
rect 15258 31226 17146 31466
rect 20212 31266 21770 31506
rect 24424 31288 26368 31528
rect 29781 31132 29983 31133
rect 30372 31132 30572 35653
rect 29781 30932 29782 31132
rect 29982 30932 30572 31132
rect 29781 30931 29983 30932
rect 11186 30678 30292 30742
rect 11016 30508 25628 30568
rect 10802 30322 21042 30382
rect 30232 30361 30292 30678
rect 30229 30360 30295 30361
rect 30229 30296 30230 30360
rect 30294 30296 30295 30360
rect 30229 30295 30295 30296
rect 10580 30132 16404 30192
rect 11428 28467 11630 28468
rect 11428 28462 11429 28467
rect 9800 28262 11429 28462
rect 1168 27556 1372 27557
rect 200 27354 1169 27556
rect 1371 27354 1372 27556
rect 200 7520 500 27354
rect 1168 27353 1372 27354
rect 200 7220 8674 7520
rect 200 1000 500 7220
rect 8374 5928 8674 7220
rect 8374 5927 9350 5928
rect 8374 5629 9051 5927
rect 9349 5629 9350 5927
rect 8374 5628 9350 5629
rect 9800 2411 10100 28262
rect 11428 28257 11429 28262
rect 11629 28257 11630 28467
rect 11428 28256 11630 28257
rect 29431 25994 29633 25995
rect 30372 25994 30572 30932
rect 29431 25794 29432 25994
rect 29632 25794 30572 25994
rect 29431 25793 29633 25794
rect 12453 4100 12727 4101
rect 12453 3828 12454 4100
rect 12726 3828 12727 4100
rect 9800 2113 9801 2411
rect 10099 2113 10100 2411
rect 9800 462 10100 2113
rect 10255 3749 10520 3750
rect 10255 3486 10256 3749
rect 10519 3486 10520 3749
rect 10255 273 10520 3486
rect 400 0 520 200
rect 4816 0 4936 200
rect 9160 120 10520 273
rect 12453 277 12727 3828
rect 30372 644 30572 25794
rect 30372 444 31412 644
rect 12453 120 13845 277
rect 31212 228 31412 444
rect 9158 0 10520 120
rect 12452 0 13846 120
rect 18064 0 18184 200
rect 22480 0 22600 200
rect 26896 0 27016 200
rect 31200 0 31432 228
use analog_mux  analog_mux_0 ~/Desktop/TinyTapeout/TinyTapeoutAnalog/tt06-programmable-thing/mag
timestamp 1713470770
transform 0 1 26232 -1 0 40002
box -240 -16 3910 4523
use analog_mux  analog_mux_1
timestamp 1713470770
transform 0 1 21506 -1 0 40004
box -240 -16 3910 4523
use analog_mux  analog_mux_2
timestamp 1713470770
transform 0 1 16856 -1 0 40006
box -240 -16 3910 4523
use analog_mux  analog_mux_3
timestamp 1713470770
transform 0 1 11908 -1 0 40022
box -240 -16 3910 4523
use analog_mux  analog_mux_4
timestamp 1713470770
transform 0 1 25722 -1 0 34848
box -240 -16 3910 4523
use analog_mux  analog_mux_5
timestamp 1713470770
transform 0 1 21102 -1 0 34826
box -240 -16 3910 4523
use analog_mux  analog_mux_6
timestamp 1713470770
transform 0 1 16522 -1 0 34786
box -240 -16 3910 4523
use analog_mux  analog_mux_7
timestamp 1713470770
transform 0 1 11886 -1 0 34804
box -240 -16 3910 4523
use analog_mux  analog_mux_8
timestamp 1713470770
transform 0 1 25772 -1 0 29704
box -240 -16 3910 4523
use inverter  inverter_0 ~/Desktop/TinyTapeout/TinyTapeoutAnalog/tt06-programmable-thing/mag
timestamp 1713454966
transform 1 0 11228 0 1 864
box -560 20 1088 6242
<< labels >>
flabel metal4 s 30974 44952 31034 45152 0 FreeSans 480 90 0 0 clk
port 0 nsew signal input
flabel metal4 s 31710 44952 31770 45152 0 FreeSans 480 90 0 0 ena
port 1 nsew signal input
flabel metal4 s 30238 44952 30298 45152 0 FreeSans 480 90 0 0 rst_n
port 2 nsew signal input
flabel metal4 s 31312 0 31432 200 0 FreeSans 960 0 0 0 ua[0]
port 3 nsew signal bidirectional
flabel metal4 s 26896 0 27016 200 0 FreeSans 960 0 0 0 ua[1]
port 4 nsew signal bidirectional
flabel metal4 s 22480 0 22600 200 0 FreeSans 960 0 0 0 ua[2]
port 5 nsew signal bidirectional
flabel metal4 s 18064 0 18184 200 0 FreeSans 960 0 0 0 ua[3]
port 6 nsew signal bidirectional
flabel metal4 s 13648 0 13768 200 0 FreeSans 960 0 0 0 ua[4]
port 7 nsew signal bidirectional
flabel metal4 s 9232 0 9352 200 0 FreeSans 960 0 0 0 ua[5]
port 8 nsew signal bidirectional
flabel metal4 s 4816 0 4936 200 0 FreeSans 960 0 0 0 ua[6]
port 9 nsew signal bidirectional
flabel metal4 s 400 0 520 200 0 FreeSans 960 0 0 0 ua[7]
port 10 nsew signal bidirectional
flabel metal4 s 29502 44952 29562 45152 0 FreeSans 480 90 0 0 ui_in[0]
port 11 nsew signal input
flabel metal4 s 28766 44952 28826 45152 0 FreeSans 480 90 0 0 ui_in[1]
port 12 nsew signal input
flabel metal4 s 28030 44952 28090 45152 0 FreeSans 480 90 0 0 ui_in[2]
port 13 nsew signal input
flabel metal4 s 27294 44952 27354 45152 0 FreeSans 480 90 0 0 ui_in[3]
port 14 nsew signal input
flabel metal4 s 26558 44952 26618 45152 0 FreeSans 480 90 0 0 ui_in[4]
port 15 nsew signal input
flabel metal4 s 25822 44952 25882 45152 0 FreeSans 480 90 0 0 ui_in[5]
port 16 nsew signal input
flabel metal4 s 25086 44952 25146 45152 0 FreeSans 480 90 0 0 ui_in[6]
port 17 nsew signal input
flabel metal4 s 24350 44952 24410 45152 0 FreeSans 480 90 0 0 ui_in[7]
port 18 nsew signal input
flabel metal4 s 23614 44952 23674 45152 0 FreeSans 480 90 0 0 uio_in[0]
port 19 nsew signal input
flabel metal4 s 22878 44952 22938 45152 0 FreeSans 480 90 0 0 uio_in[1]
port 20 nsew signal input
flabel metal4 s 22142 44952 22202 45152 0 FreeSans 480 90 0 0 uio_in[2]
port 21 nsew signal input
flabel metal4 s 21406 44952 21466 45152 0 FreeSans 480 90 0 0 uio_in[3]
port 22 nsew signal input
flabel metal4 s 20670 44952 20730 45152 0 FreeSans 480 90 0 0 uio_in[4]
port 23 nsew signal input
flabel metal4 s 19934 44952 19994 45152 0 FreeSans 480 90 0 0 uio_in[5]
port 24 nsew signal input
flabel metal4 s 19198 44952 19258 45152 0 FreeSans 480 90 0 0 uio_in[6]
port 25 nsew signal input
flabel metal4 s 18462 44952 18522 45152 0 FreeSans 480 90 0 0 uio_in[7]
port 26 nsew signal input
flabel metal4 s 5950 44952 6010 45152 0 FreeSans 480 90 0 0 uio_oe[0]
port 27 nsew signal output
flabel metal4 s 5214 44952 5274 45152 0 FreeSans 480 90 0 0 uio_oe[1]
port 28 nsew signal output
flabel metal4 s 4478 44952 4538 45152 0 FreeSans 480 90 0 0 uio_oe[2]
port 29 nsew signal output
flabel metal4 s 3742 44952 3802 45152 0 FreeSans 480 90 0 0 uio_oe[3]
port 30 nsew signal output
flabel metal4 s 3006 44952 3066 45152 0 FreeSans 480 90 0 0 uio_oe[4]
port 31 nsew signal output
flabel metal4 s 2270 44952 2330 45152 0 FreeSans 480 90 0 0 uio_oe[5]
port 32 nsew signal output
flabel metal4 s 1534 44952 1594 45152 0 FreeSans 480 90 0 0 uio_oe[6]
port 33 nsew signal output
flabel metal4 s 798 44952 858 45152 0 FreeSans 480 90 0 0 uio_oe[7]
port 34 nsew signal output
flabel metal4 s 11838 44952 11898 45152 0 FreeSans 480 90 0 0 uio_out[0]
port 35 nsew signal output
flabel metal4 s 11102 44952 11162 45152 0 FreeSans 480 90 0 0 uio_out[1]
port 36 nsew signal output
flabel metal4 s 10366 44952 10426 45152 0 FreeSans 480 90 0 0 uio_out[2]
port 37 nsew signal output
flabel metal4 s 9630 44952 9690 45152 0 FreeSans 480 90 0 0 uio_out[3]
port 38 nsew signal output
flabel metal4 s 8894 44952 8954 45152 0 FreeSans 480 90 0 0 uio_out[4]
port 39 nsew signal output
flabel metal4 s 8158 44952 8218 45152 0 FreeSans 480 90 0 0 uio_out[5]
port 40 nsew signal output
flabel metal4 s 7422 44952 7482 45152 0 FreeSans 480 90 0 0 uio_out[6]
port 41 nsew signal output
flabel metal4 s 6686 44952 6746 45152 0 FreeSans 480 90 0 0 uio_out[7]
port 42 nsew signal output
flabel metal4 s 17726 44952 17786 45152 0 FreeSans 480 90 0 0 uo_out[0]
port 43 nsew signal output
flabel metal4 s 16990 44952 17050 45152 0 FreeSans 480 90 0 0 uo_out[1]
port 44 nsew signal output
flabel metal4 s 16254 44952 16314 45152 0 FreeSans 480 90 0 0 uo_out[2]
port 45 nsew signal output
flabel metal4 s 15518 44952 15578 45152 0 FreeSans 480 90 0 0 uo_out[3]
port 46 nsew signal output
flabel metal4 s 14782 44952 14842 45152 0 FreeSans 480 90 0 0 uo_out[4]
port 47 nsew signal output
flabel metal4 s 14046 44952 14106 45152 0 FreeSans 480 90 0 0 uo_out[5]
port 48 nsew signal output
flabel metal4 s 13310 44952 13370 45152 0 FreeSans 480 90 0 0 uo_out[6]
port 49 nsew signal output
flabel metal4 s 12574 44952 12634 45152 0 FreeSans 480 90 0 0 uo_out[7]
port 50 nsew signal output
flabel metal4 200 1000 500 44152 1 FreeSans 2 0 0 0 VPWR
port 51 nsew power bidirectional
flabel metal4 9800 1000 10100 44152 1 FreeSans 2 0 0 0 VGND
port 52 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 32200 45152
<< end >>
