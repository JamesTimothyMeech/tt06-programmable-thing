VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO tt_um_JamesTimothyMeech_inverter
  CLASS BLOCK ;
  FOREIGN tt_um_JamesTimothyMeech_inverter ;
  ORIGIN 0.000 0.000 ;
  SIZE 161.000 BY 225.760 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 154.870 224.760 155.170 225.760 ;
    END
  END clk
  PIN ena
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 158.550 224.760 158.850 225.760 ;
    END
  END ena
  PIN rst_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 151.190 224.760 151.490 225.760 ;
    END
  END rst_n
  PIN ua[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 156.560 0.000 157.160 1.000 ;
    END
  END ua[0]
  PIN ua[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 134.480 0.000 135.080 1.000 ;
    END
  END ua[1]
  PIN ua[2]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 112.400 0.000 113.000 1.000 ;
    END
  END ua[2]
  PIN ua[3]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 90.320 0.000 90.920 1.000 ;
    END
  END ua[3]
  PIN ua[4]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 5.800000 ;
    PORT
      LAYER met4 ;
        RECT 68.240 0.000 68.840 1.000 ;
    END
  END ua[4]
  PIN ua[5]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 20.000000 ;
    PORT
      LAYER met4 ;
        RECT 46.160 0.000 46.760 1.000 ;
    END
  END ua[5]
  PIN ua[6]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 24.080 0.000 24.680 1.000 ;
    END
  END ua[6]
  PIN ua[7]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 2.000 0.000 2.600 1.000 ;
    END
  END ua[7]
  PIN ui_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 147.510 224.760 147.810 225.760 ;
    END
  END ui_in[0]
  PIN ui_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 143.830 224.760 144.130 225.760 ;
    END
  END ui_in[1]
  PIN ui_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 140.150 224.760 140.450 225.760 ;
    END
  END ui_in[2]
  PIN ui_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 136.470 224.760 136.770 225.760 ;
    END
  END ui_in[3]
  PIN ui_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 132.790 224.760 133.090 225.760 ;
    END
  END ui_in[4]
  PIN ui_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 129.110 224.760 129.410 225.760 ;
    END
  END ui_in[5]
  PIN ui_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 125.430 224.760 125.730 225.760 ;
    END
  END ui_in[6]
  PIN ui_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 121.750 224.760 122.050 225.760 ;
    END
  END ui_in[7]
  PIN uio_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 118.070 224.760 118.370 225.760 ;
    END
  END uio_in[0]
  PIN uio_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 114.390 224.760 114.690 225.760 ;
    END
  END uio_in[1]
  PIN uio_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 110.710 224.760 111.010 225.760 ;
    END
  END uio_in[2]
  PIN uio_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 107.030 224.760 107.330 225.760 ;
    END
  END uio_in[3]
  PIN uio_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 103.350 224.760 103.650 225.760 ;
    END
  END uio_in[4]
  PIN uio_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 99.670 224.760 99.970 225.760 ;
    END
  END uio_in[5]
  PIN uio_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 95.990 224.760 96.290 225.760 ;
    END
  END uio_in[6]
  PIN uio_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 92.310 224.760 92.610 225.760 ;
    END
  END uio_in[7]
  PIN uio_oe[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 29.750 224.760 30.050 225.760 ;
    END
  END uio_oe[0]
  PIN uio_oe[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 26.070 224.760 26.370 225.760 ;
    END
  END uio_oe[1]
  PIN uio_oe[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 22.390 224.760 22.690 225.760 ;
    END
  END uio_oe[2]
  PIN uio_oe[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 18.710 224.760 19.010 225.760 ;
    END
  END uio_oe[3]
  PIN uio_oe[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 15.030 224.760 15.330 225.760 ;
    END
  END uio_oe[4]
  PIN uio_oe[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 11.350 224.760 11.650 225.760 ;
    END
  END uio_oe[5]
  PIN uio_oe[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 7.670 224.760 7.970 225.760 ;
    END
  END uio_oe[6]
  PIN uio_oe[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 3.990 224.760 4.290 225.760 ;
    END
  END uio_oe[7]
  PIN uio_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 59.190 224.760 59.490 225.760 ;
    END
  END uio_out[0]
  PIN uio_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 55.510 224.760 55.810 225.760 ;
    END
  END uio_out[1]
  PIN uio_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 51.830 224.760 52.130 225.760 ;
    END
  END uio_out[2]
  PIN uio_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 48.150 224.760 48.450 225.760 ;
    END
  END uio_out[3]
  PIN uio_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 44.470 224.760 44.770 225.760 ;
    END
  END uio_out[4]
  PIN uio_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 40.790 224.760 41.090 225.760 ;
    END
  END uio_out[5]
  PIN uio_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 37.110 224.760 37.410 225.760 ;
    END
  END uio_out[6]
  PIN uio_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 33.430 224.760 33.730 225.760 ;
    END
  END uio_out[7]
  PIN uo_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 88.630 224.760 88.930 225.760 ;
    END
  END uo_out[0]
  PIN uo_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 84.950 224.760 85.250 225.760 ;
    END
  END uo_out[1]
  PIN uo_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 81.270 224.760 81.570 225.760 ;
    END
  END uo_out[2]
  PIN uo_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 77.590 224.760 77.890 225.760 ;
    END
  END uo_out[3]
  PIN uo_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 73.910 224.760 74.210 225.760 ;
    END
  END uo_out[4]
  PIN uo_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 70.230 224.760 70.530 225.760 ;
    END
  END uo_out[5]
  PIN uo_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 66.550 224.760 66.850 225.760 ;
    END
  END uo_out[6]
  PIN uo_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 62.870 224.760 63.170 225.760 ;
    END
  END uo_out[7]
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1.000 5.000 2.500 220.760 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 49.000 5.000 50.500 220.760 ;
    END
  END VGND
  OBS
      LAYER nwell ;
        RECT 57.550 22.720 60.510 34.910 ;
      LAYER pwell ;
        RECT 57.500 16.280 60.460 17.430 ;
        RECT 57.500 6.480 60.520 16.280 ;
        RECT 57.500 5.330 60.460 6.480 ;
      LAYER li1 ;
        RECT 57.730 34.560 60.330 34.730 ;
        RECT 57.730 33.600 57.900 34.560 ;
        RECT 58.530 34.050 59.530 34.220 ;
        RECT 57.730 23.990 57.910 33.600 ;
        RECT 57.730 23.070 57.900 23.990 ;
        RECT 58.300 23.795 58.470 33.835 ;
        RECT 59.590 23.795 59.760 33.835 ;
        RECT 58.530 23.410 59.530 23.580 ;
        RECT 60.160 23.070 60.330 34.560 ;
        RECT 57.730 22.900 60.330 23.070 ;
        RECT 57.680 17.080 60.280 17.250 ;
        RECT 57.680 5.680 57.850 17.080 ;
        RECT 58.480 16.570 59.480 16.740 ;
        RECT 58.250 6.360 58.420 16.400 ;
        RECT 59.540 6.360 59.710 16.400 ;
        RECT 58.480 6.020 59.480 6.190 ;
        RECT 60.110 5.680 60.280 17.080 ;
        RECT 57.680 5.510 60.280 5.680 ;
      LAYER mcon ;
        RECT 58.210 34.560 59.850 34.730 ;
        RECT 58.610 34.050 59.450 34.220 ;
        RECT 57.740 23.990 57.910 33.600 ;
        RECT 58.300 23.875 58.470 33.755 ;
        RECT 59.590 23.875 59.760 33.755 ;
        RECT 58.610 23.410 59.450 23.580 ;
        RECT 58.560 16.570 59.400 16.740 ;
        RECT 57.680 6.630 57.850 16.130 ;
        RECT 58.250 6.440 58.420 16.320 ;
        RECT 59.540 6.440 59.710 16.320 ;
        RECT 58.560 6.020 59.400 6.190 ;
        RECT 58.160 5.510 59.800 5.680 ;
      LAYER met1 ;
        RECT 43.900 36.070 45.400 37.630 ;
        RECT 44.125 35.490 45.135 36.070 ;
        RECT 55.080 35.490 55.720 35.510 ;
        RECT 56.285 35.490 56.925 35.500 ;
        RECT 44.125 34.540 60.520 35.490 ;
        RECT 44.125 34.490 60.500 34.540 ;
        RECT 44.125 34.480 57.340 34.490 ;
        RECT 54.610 34.470 56.900 34.480 ;
        RECT 58.550 34.220 59.510 34.250 ;
        RECT 53.345 34.050 59.510 34.220 ;
        RECT 53.345 23.580 53.750 34.050 ;
        RECT 58.550 34.020 59.510 34.050 ;
        RECT 58.270 33.760 58.500 33.815 ;
        RECT 54.050 23.870 58.500 33.760 ;
        RECT 58.270 23.815 58.500 23.870 ;
        RECT 59.560 33.760 59.790 33.815 ;
        RECT 59.560 23.870 61.580 33.760 ;
        RECT 59.560 23.815 59.790 23.870 ;
        RECT 58.550 23.580 59.510 23.610 ;
        RECT 53.345 23.410 59.510 23.580 ;
        RECT 53.345 20.510 54.345 23.410 ;
        RECT 58.550 23.380 59.510 23.410 ;
        RECT 60.590 20.535 61.580 23.870 ;
        RECT 53.245 19.125 54.570 20.510 ;
        RECT 53.345 16.740 54.345 19.125 ;
        RECT 60.395 19.105 61.765 20.535 ;
        RECT 60.590 18.395 61.580 19.105 ;
        RECT 58.500 16.740 59.460 16.770 ;
        RECT 53.345 16.570 59.480 16.740 ;
        RECT 53.345 6.190 53.750 16.570 ;
        RECT 58.500 16.540 59.460 16.570 ;
        RECT 58.220 16.280 58.450 16.380 ;
        RECT 54.030 6.480 58.450 16.280 ;
        RECT 54.595 6.455 57.050 6.480 ;
        RECT 54.625 6.415 57.020 6.455 ;
        RECT 58.220 6.380 58.450 6.480 ;
        RECT 59.510 16.280 59.740 16.380 ;
        RECT 60.610 16.280 61.575 18.395 ;
        RECT 59.510 6.480 61.575 16.280 ;
        RECT 59.510 6.380 59.740 6.480 ;
        RECT 58.500 6.190 59.460 6.220 ;
        RECT 53.345 6.015 59.460 6.190 ;
        RECT 53.345 6.010 53.750 6.015 ;
        RECT 58.500 5.990 59.460 6.015 ;
        RECT 54.600 5.820 55.185 5.850 ;
        RECT 55.685 5.820 57.030 5.850 ;
        RECT 54.600 5.800 57.060 5.820 ;
        RECT 48.980 4.800 60.460 5.800 ;
        RECT 49.000 4.790 60.460 4.800 ;
        RECT 49.000 3.630 60.440 4.790 ;
        RECT 49.000 3.600 50.500 3.630 ;
      LAYER via ;
        RECT 43.900 36.100 45.400 37.600 ;
        RECT 55.110 35.490 55.690 35.510 ;
        RECT 56.315 35.490 56.895 35.500 ;
        RECT 54.610 34.920 56.895 35.490 ;
        RECT 54.610 34.490 56.870 34.920 ;
        RECT 54.610 24.390 56.895 33.710 ;
        RECT 53.245 19.155 54.570 20.480 ;
        RECT 60.395 19.135 61.765 20.505 ;
        RECT 54.625 6.455 57.020 15.765 ;
        RECT 54.600 5.375 57.030 5.820 ;
        RECT 54.600 4.790 57.040 5.375 ;
        RECT 55.080 4.760 56.640 4.790 ;
      LAYER met2 ;
        RECT 43.925 37.600 45.375 37.620 ;
        RECT 43.870 36.100 45.430 37.600 ;
        RECT 43.925 36.080 45.375 36.100 ;
        RECT 55.110 35.520 55.690 35.540 ;
        RECT 56.315 35.520 56.895 35.530 ;
        RECT 54.610 24.360 56.895 35.520 ;
        RECT 62.290 20.505 63.610 20.525 ;
        RECT 51.300 20.480 52.575 20.500 ;
        RECT 51.275 19.155 54.600 20.480 ;
        RECT 51.300 19.135 52.575 19.155 ;
        RECT 60.365 19.135 63.635 20.505 ;
        RECT 62.290 19.115 63.610 19.135 ;
        RECT 54.625 11.135 57.020 15.805 ;
        RECT 49.000 6.735 50.500 6.760 ;
        RECT 48.980 5.285 50.520 6.735 ;
        RECT 54.595 6.455 57.050 11.135 ;
        RECT 54.600 5.820 57.030 6.455 ;
        RECT 54.570 5.375 57.060 5.820 ;
        RECT 49.000 5.130 50.500 5.285 ;
        RECT 54.570 5.235 57.070 5.375 ;
        RECT 48.970 3.630 50.530 5.130 ;
        RECT 54.600 4.790 57.070 5.235 ;
        RECT 54.600 4.760 57.040 4.790 ;
        RECT 55.080 4.750 55.665 4.760 ;
      LAYER via2 ;
        RECT 43.925 36.125 45.375 37.575 ;
        RECT 51.300 19.180 52.575 20.455 ;
        RECT 62.290 19.160 63.610 20.480 ;
        RECT 49.025 5.285 50.475 6.735 ;
      LAYER met3 ;
        RECT 43.905 37.600 45.395 37.625 ;
        RECT 43.900 36.100 45.400 37.600 ;
        RECT 43.905 36.075 45.395 36.100 ;
        RECT 62.265 20.500 63.635 20.505 ;
        RECT 51.275 20.475 52.600 20.480 ;
        RECT 51.250 19.160 52.625 20.475 ;
        RECT 51.275 19.155 52.600 19.160 ;
        RECT 62.240 19.140 63.660 20.500 ;
        RECT 62.265 19.135 63.635 19.140 ;
        RECT 49.000 6.755 50.500 6.760 ;
        RECT 48.975 5.265 50.525 6.755 ;
        RECT 49.000 5.260 50.500 5.265 ;
      LAYER via3 ;
        RECT 43.905 36.105 45.395 37.595 ;
        RECT 51.280 19.160 52.595 20.475 ;
        RECT 62.270 19.140 63.630 20.500 ;
        RECT 49.005 5.265 50.495 6.755 ;
      LAYER met4 ;
        RECT 3.990 223.390 4.290 224.760 ;
        RECT 7.670 223.390 7.970 224.760 ;
        RECT 11.350 223.390 11.650 224.760 ;
        RECT 15.030 223.390 15.330 224.760 ;
        RECT 18.710 223.390 19.010 224.760 ;
        RECT 22.390 223.390 22.690 224.760 ;
        RECT 26.070 223.390 26.370 224.760 ;
        RECT 29.750 223.390 30.050 224.760 ;
        RECT 33.430 223.390 33.730 224.760 ;
        RECT 37.110 223.390 37.410 224.760 ;
        RECT 40.790 223.390 41.090 224.760 ;
        RECT 44.470 223.390 44.770 224.760 ;
        RECT 48.150 223.390 48.450 224.760 ;
        RECT 51.830 223.390 52.130 224.760 ;
        RECT 55.510 223.390 55.810 224.760 ;
        RECT 59.190 223.390 59.490 224.760 ;
        RECT 62.870 223.390 63.170 224.760 ;
        RECT 66.550 223.390 66.850 224.760 ;
        RECT 70.230 223.390 70.530 224.760 ;
        RECT 73.910 223.390 74.210 224.760 ;
        RECT 77.590 223.390 77.890 224.760 ;
        RECT 81.270 223.390 81.570 224.760 ;
        RECT 84.950 223.390 85.250 224.760 ;
        RECT 88.630 223.390 88.930 224.760 ;
        RECT 3.385 222.320 89.730 223.390 ;
        RECT 2.500 36.100 45.400 37.600 ;
        RECT 51.275 1.365 52.600 20.480 ;
        RECT 45.800 1.000 52.600 1.365 ;
        RECT 45.800 0.040 46.160 1.000 ;
        RECT 46.760 0.040 52.600 1.000 ;
        RECT 62.265 1.385 63.635 20.505 ;
        RECT 62.265 1.000 69.225 1.385 ;
        RECT 62.265 0.015 68.240 1.000 ;
        RECT 68.840 0.015 69.225 1.000 ;
  END
END tt_um_JamesTimothyMeech_inverter
END LIBRARY

